library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NCO_ILA is
    port (
        clk_i: in std_logic;
        rst_i: in std_logic
    );
end entity NCO_ILA;

architecture NCO_ILA_arch of NCO_ILA is
        -- declarations

component NCO is
    port (
        clk_i: in std_logic;
        rst_i: in std_logic;
        pha_i: in std_logic_vector(15 downto 0);
        q_o:   out std_logic_vector(11 downto 0)
    );
end component NCO;

COMPONENT ila_0

PORT (
	clk : IN STD_LOGIC;
	probe0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0)
);
END COMPONENT  ;

COMPONENT vio_0
  PORT (
    clk : IN STD_LOGIC;
    probe_out0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

    type sin_lut_type is array (0 to 4095) of std_logic_vector(11 downto 0);
    constant sin_lut: sin_lut_type := ( 
        0 => "011111111111",
        1 => "100000000010",
        2 => "100000000101",
        3 => "100000001000",
        4 => "100000001100",
        5 => "100000001111",
        6 => "100000010010",
        7 => "100000010101",
        8 => "100000011000",
        9 => "100000011011",
        10 => "100000011110",
        11 => "100000100010",
        12 => "100000100101",
        13 => "100000101000",
        14 => "100000101011",
        15 => "100000101110",
        16 => "100000110001",
        17 => "100000110100",
        18 => "100000111000",
        19 => "100000111011",
        20 => "100000111110",
        21 => "100001000001",
        22 => "100001000100",
        23 => "100001000111",
        24 => "100001001010",
        25 => "100001001110",
        26 => "100001010001",
        27 => "100001010100",
        28 => "100001010111",
        29 => "100001011010",
        30 => "100001011101",
        31 => "100001100000",
        32 => "100001100011",
        33 => "100001100111",
        34 => "100001101010",
        35 => "100001101101",
        36 => "100001110000",
        37 => "100001110011",
        38 => "100001110110",
        39 => "100001111001",
        40 => "100001111101",
        41 => "100010000000",
        42 => "100010000011",
        43 => "100010000110",
        44 => "100010001001",
        45 => "100010001100",
        46 => "100010001111",
        47 => "100010010010",
        48 => "100010010110",
        49 => "100010011001",
        50 => "100010011100",
        51 => "100010011111",
        52 => "100010100010",
        53 => "100010100101",
        54 => "100010101000",
        55 => "100010101100",
        56 => "100010101111",
        57 => "100010110010",
        58 => "100010110101",
        59 => "100010111000",
        60 => "100010111011",
        61 => "100010111110",
        62 => "100011000001",
        63 => "100011000101",
        64 => "100011001000",
        65 => "100011001011",
        66 => "100011001110",
        67 => "100011010001",
        68 => "100011010100",
        69 => "100011010111",
        70 => "100011011010",
        71 => "100011011110",
        72 => "100011100001",
        73 => "100011100100",
        74 => "100011100111",
        75 => "100011101010",
        76 => "100011101101",
        77 => "100011110000",
        78 => "100011110011",
        79 => "100011110111",
        80 => "100011111010",
        81 => "100011111101",
        82 => "100100000000",
        83 => "100100000011",
        84 => "100100000110",
        85 => "100100001001",
        86 => "100100001100",
        87 => "100100001111",
        88 => "100100010011",
        89 => "100100010110",
        90 => "100100011001",
        91 => "100100011100",
        92 => "100100011111",
        93 => "100100100010",
        94 => "100100100101",
        95 => "100100101000",
        96 => "100100101011",
        97 => "100100101111",
        98 => "100100110010",
        99 => "100100110101",
        100 => "100100111000",
        101 => "100100111011",
        102 => "100100111110",
        103 => "100101000001",
        104 => "100101000100",
        105 => "100101000111",
        106 => "100101001010",
        107 => "100101001110",
        108 => "100101010001",
        109 => "100101010100",
        110 => "100101010111",
        111 => "100101011010",
        112 => "100101011101",
        113 => "100101100000",
        114 => "100101100011",
        115 => "100101100110",
        116 => "100101101001",
        117 => "100101101101",
        118 => "100101110000",
        119 => "100101110011",
        120 => "100101110110",
        121 => "100101111001",
        122 => "100101111100",
        123 => "100101111111",
        124 => "100110000010",
        125 => "100110000101",
        126 => "100110001000",
        127 => "100110001011",
        128 => "100110001110",
        129 => "100110010010",
        130 => "100110010101",
        131 => "100110011000",
        132 => "100110011011",
        133 => "100110011110",
        134 => "100110100001",
        135 => "100110100100",
        136 => "100110100111",
        137 => "100110101010",
        138 => "100110101101",
        139 => "100110110000",
        140 => "100110110011",
        141 => "100110110110",
        142 => "100110111001",
        143 => "100110111101",
        144 => "100111000000",
        145 => "100111000011",
        146 => "100111000110",
        147 => "100111001001",
        148 => "100111001100",
        149 => "100111001111",
        150 => "100111010010",
        151 => "100111010101",
        152 => "100111011000",
        153 => "100111011011",
        154 => "100111011110",
        155 => "100111100001",
        156 => "100111100100",
        157 => "100111100111",
        158 => "100111101010",
        159 => "100111101101",
        160 => "100111110001",
        161 => "100111110100",
        162 => "100111110111",
        163 => "100111111010",
        164 => "100111111101",
        165 => "101000000000",
        166 => "101000000011",
        167 => "101000000110",
        168 => "101000001001",
        169 => "101000001100",
        170 => "101000001111",
        171 => "101000010010",
        172 => "101000010101",
        173 => "101000011000",
        174 => "101000011011",
        175 => "101000011110",
        176 => "101000100001",
        177 => "101000100100",
        178 => "101000100111",
        179 => "101000101010",
        180 => "101000101101",
        181 => "101000110000",
        182 => "101000110011",
        183 => "101000110110",
        184 => "101000111001",
        185 => "101000111100",
        186 => "101000111111",
        187 => "101001000010",
        188 => "101001000101",
        189 => "101001001000",
        190 => "101001001011",
        191 => "101001001110",
        192 => "101001010001",
        193 => "101001010100",
        194 => "101001010111",
        195 => "101001011010",
        196 => "101001011101",
        197 => "101001100000",
        198 => "101001100011",
        199 => "101001100110",
        200 => "101001101001",
        201 => "101001101100",
        202 => "101001101111",
        203 => "101001110010",
        204 => "101001110101",
        205 => "101001111000",
        206 => "101001111011",
        207 => "101001111110",
        208 => "101010000001",
        209 => "101010000100",
        210 => "101010000111",
        211 => "101010001010",
        212 => "101010001101",
        213 => "101010010000",
        214 => "101010010011",
        215 => "101010010110",
        216 => "101010011001",
        217 => "101010011100",
        218 => "101010011111",
        219 => "101010100010",
        220 => "101010100101",
        221 => "101010101000",
        222 => "101010101011",
        223 => "101010101110",
        224 => "101010110001",
        225 => "101010110100",
        226 => "101010110111",
        227 => "101010111010",
        228 => "101010111101",
        229 => "101011000000",
        230 => "101011000010",
        231 => "101011000101",
        232 => "101011001000",
        233 => "101011001011",
        234 => "101011001110",
        235 => "101011010001",
        236 => "101011010100",
        237 => "101011010111",
        238 => "101011011010",
        239 => "101011011101",
        240 => "101011100000",
        241 => "101011100011",
        242 => "101011100110",
        243 => "101011101001",
        244 => "101011101100",
        245 => "101011101111",
        246 => "101011110001",
        247 => "101011110100",
        248 => "101011110111",
        249 => "101011111010",
        250 => "101011111101",
        251 => "101100000000",
        252 => "101100000011",
        253 => "101100000110",
        254 => "101100001001",
        255 => "101100001100",
        256 => "101100001111",
        257 => "101100010001",
        258 => "101100010100",
        259 => "101100010111",
        260 => "101100011010",
        261 => "101100011101",
        262 => "101100100000",
        263 => "101100100011",
        264 => "101100100110",
        265 => "101100101001",
        266 => "101100101011",
        267 => "101100101110",
        268 => "101100110001",
        269 => "101100110100",
        270 => "101100110111",
        271 => "101100111010",
        272 => "101100111101",
        273 => "101101000000",
        274 => "101101000010",
        275 => "101101000101",
        276 => "101101001000",
        277 => "101101001011",
        278 => "101101001110",
        279 => "101101010001",
        280 => "101101010100",
        281 => "101101010110",
        282 => "101101011001",
        283 => "101101011100",
        284 => "101101011111",
        285 => "101101100010",
        286 => "101101100101",
        287 => "101101101000",
        288 => "101101101010",
        289 => "101101101101",
        290 => "101101110000",
        291 => "101101110011",
        292 => "101101110110",
        293 => "101101111001",
        294 => "101101111011",
        295 => "101101111110",
        296 => "101110000001",
        297 => "101110000100",
        298 => "101110000111",
        299 => "101110001010",
        300 => "101110001100",
        301 => "101110001111",
        302 => "101110010010",
        303 => "101110010101",
        304 => "101110011000",
        305 => "101110011010",
        306 => "101110011101",
        307 => "101110100000",
        308 => "101110100011",
        309 => "101110100110",
        310 => "101110101000",
        311 => "101110101011",
        312 => "101110101110",
        313 => "101110110001",
        314 => "101110110100",
        315 => "101110110110",
        316 => "101110111001",
        317 => "101110111100",
        318 => "101110111111",
        319 => "101111000001",
        320 => "101111000100",
        321 => "101111000111",
        322 => "101111001010",
        323 => "101111001100",
        324 => "101111001111",
        325 => "101111010010",
        326 => "101111010101",
        327 => "101111011000",
        328 => "101111011010",
        329 => "101111011101",
        330 => "101111100000",
        331 => "101111100011",
        332 => "101111100101",
        333 => "101111101000",
        334 => "101111101011",
        335 => "101111101101",
        336 => "101111110000",
        337 => "101111110011",
        338 => "101111110110",
        339 => "101111111000",
        340 => "101111111011",
        341 => "101111111110",
        342 => "110000000001",
        343 => "110000000011",
        344 => "110000000110",
        345 => "110000001001",
        346 => "110000001011",
        347 => "110000001110",
        348 => "110000010001",
        349 => "110000010100",
        350 => "110000010110",
        351 => "110000011001",
        352 => "110000011100",
        353 => "110000011110",
        354 => "110000100001",
        355 => "110000100100",
        356 => "110000100110",
        357 => "110000101001",
        358 => "110000101100",
        359 => "110000101110",
        360 => "110000110001",
        361 => "110000110100",
        362 => "110000110110",
        363 => "110000111001",
        364 => "110000111100",
        365 => "110000111110",
        366 => "110001000001",
        367 => "110001000100",
        368 => "110001000110",
        369 => "110001001001",
        370 => "110001001100",
        371 => "110001001110",
        372 => "110001010001",
        373 => "110001010100",
        374 => "110001010110",
        375 => "110001011001",
        376 => "110001011100",
        377 => "110001011110",
        378 => "110001100001",
        379 => "110001100011",
        380 => "110001100110",
        381 => "110001101001",
        382 => "110001101011",
        383 => "110001101110",
        384 => "110001110001",
        385 => "110001110011",
        386 => "110001110110",
        387 => "110001111000",
        388 => "110001111011",
        389 => "110001111110",
        390 => "110010000000",
        391 => "110010000011",
        392 => "110010000101",
        393 => "110010001000",
        394 => "110010001011",
        395 => "110010001101",
        396 => "110010010000",
        397 => "110010010010",
        398 => "110010010101",
        399 => "110010010111",
        400 => "110010011010",
        401 => "110010011101",
        402 => "110010011111",
        403 => "110010100010",
        404 => "110010100100",
        405 => "110010100111",
        406 => "110010101001",
        407 => "110010101100",
        408 => "110010101110",
        409 => "110010110001",
        410 => "110010110100",
        411 => "110010110110",
        412 => "110010111001",
        413 => "110010111011",
        414 => "110010111110",
        415 => "110011000000",
        416 => "110011000011",
        417 => "110011000101",
        418 => "110011001000",
        419 => "110011001010",
        420 => "110011001101",
        421 => "110011001111",
        422 => "110011010010",
        423 => "110011010100",
        424 => "110011010111",
        425 => "110011011001",
        426 => "110011011100",
        427 => "110011011110",
        428 => "110011100001",
        429 => "110011100011",
        430 => "110011100110",
        431 => "110011101000",
        432 => "110011101011",
        433 => "110011101101",
        434 => "110011110000",
        435 => "110011110010",
        436 => "110011110101",
        437 => "110011110111",
        438 => "110011111001",
        439 => "110011111100",
        440 => "110011111110",
        441 => "110100000001",
        442 => "110100000011",
        443 => "110100000110",
        444 => "110100001000",
        445 => "110100001011",
        446 => "110100001101",
        447 => "110100001111",
        448 => "110100010010",
        449 => "110100010100",
        450 => "110100010111",
        451 => "110100011001",
        452 => "110100011100",
        453 => "110100011110",
        454 => "110100100000",
        455 => "110100100011",
        456 => "110100100101",
        457 => "110100101000",
        458 => "110100101010",
        459 => "110100101100",
        460 => "110100101111",
        461 => "110100110001",
        462 => "110100110100",
        463 => "110100110110",
        464 => "110100111000",
        465 => "110100111011",
        466 => "110100111101",
        467 => "110100111111",
        468 => "110101000010",
        469 => "110101000100",
        470 => "110101000111",
        471 => "110101001001",
        472 => "110101001011",
        473 => "110101001110",
        474 => "110101010000",
        475 => "110101010010",
        476 => "110101010101",
        477 => "110101010111",
        478 => "110101011001",
        479 => "110101011100",
        480 => "110101011110",
        481 => "110101100000",
        482 => "110101100011",
        483 => "110101100101",
        484 => "110101100111",
        485 => "110101101010",
        486 => "110101101100",
        487 => "110101101110",
        488 => "110101110001",
        489 => "110101110011",
        490 => "110101110101",
        491 => "110101110111",
        492 => "110101111010",
        493 => "110101111100",
        494 => "110101111110",
        495 => "110110000001",
        496 => "110110000011",
        497 => "110110000101",
        498 => "110110000111",
        499 => "110110001010",
        500 => "110110001100",
        501 => "110110001110",
        502 => "110110010000",
        503 => "110110010011",
        504 => "110110010101",
        505 => "110110010111",
        506 => "110110011001",
        507 => "110110011100",
        508 => "110110011110",
        509 => "110110100000",
        510 => "110110100010",
        511 => "110110100101",
        512 => "110110100111",
        513 => "110110101001",
        514 => "110110101011",
        515 => "110110101101",
        516 => "110110110000",
        517 => "110110110010",
        518 => "110110110100",
        519 => "110110110110",
        520 => "110110111000",
        521 => "110110111011",
        522 => "110110111101",
        523 => "110110111111",
        524 => "110111000001",
        525 => "110111000011",
        526 => "110111000110",
        527 => "110111001000",
        528 => "110111001010",
        529 => "110111001100",
        530 => "110111001110",
        531 => "110111010000",
        532 => "110111010011",
        533 => "110111010101",
        534 => "110111010111",
        535 => "110111011001",
        536 => "110111011011",
        537 => "110111011101",
        538 => "110111011111",
        539 => "110111100010",
        540 => "110111100100",
        541 => "110111100110",
        542 => "110111101000",
        543 => "110111101010",
        544 => "110111101100",
        545 => "110111101110",
        546 => "110111110000",
        547 => "110111110010",
        548 => "110111110101",
        549 => "110111110111",
        550 => "110111111001",
        551 => "110111111011",
        552 => "110111111101",
        553 => "110111111111",
        554 => "111000000001",
        555 => "111000000011",
        556 => "111000000101",
        557 => "111000000111",
        558 => "111000001001",
        559 => "111000001011",
        560 => "111000001101",
        561 => "111000001111",
        562 => "111000010001",
        563 => "111000010100",
        564 => "111000010110",
        565 => "111000011000",
        566 => "111000011010",
        567 => "111000011100",
        568 => "111000011110",
        569 => "111000100000",
        570 => "111000100010",
        571 => "111000100100",
        572 => "111000100110",
        573 => "111000101000",
        574 => "111000101010",
        575 => "111000101100",
        576 => "111000101110",
        577 => "111000110000",
        578 => "111000110010",
        579 => "111000110100",
        580 => "111000110110",
        581 => "111000111000",
        582 => "111000111010",
        583 => "111000111100",
        584 => "111000111110",
        585 => "111001000000",
        586 => "111001000001",
        587 => "111001000011",
        588 => "111001000101",
        589 => "111001000111",
        590 => "111001001001",
        591 => "111001001011",
        592 => "111001001101",
        593 => "111001001111",
        594 => "111001010001",
        595 => "111001010011",
        596 => "111001010101",
        597 => "111001010111",
        598 => "111001011001",
        599 => "111001011011",
        600 => "111001011100",
        601 => "111001011110",
        602 => "111001100000",
        603 => "111001100010",
        604 => "111001100100",
        605 => "111001100110",
        606 => "111001101000",
        607 => "111001101010",
        608 => "111001101100",
        609 => "111001101101",
        610 => "111001101111",
        611 => "111001110001",
        612 => "111001110011",
        613 => "111001110101",
        614 => "111001110111",
        615 => "111001111001",
        616 => "111001111010",
        617 => "111001111100",
        618 => "111001111110",
        619 => "111010000000",
        620 => "111010000010",
        621 => "111010000100",
        622 => "111010000101",
        623 => "111010000111",
        624 => "111010001001",
        625 => "111010001011",
        626 => "111010001101",
        627 => "111010001110",
        628 => "111010010000",
        629 => "111010010010",
        630 => "111010010100",
        631 => "111010010110",
        632 => "111010010111",
        633 => "111010011001",
        634 => "111010011011",
        635 => "111010011101",
        636 => "111010011110",
        637 => "111010100000",
        638 => "111010100010",
        639 => "111010100100",
        640 => "111010100101",
        641 => "111010100111",
        642 => "111010101001",
        643 => "111010101011",
        644 => "111010101100",
        645 => "111010101110",
        646 => "111010110000",
        647 => "111010110010",
        648 => "111010110011",
        649 => "111010110101",
        650 => "111010110111",
        651 => "111010111000",
        652 => "111010111010",
        653 => "111010111100",
        654 => "111010111101",
        655 => "111010111111",
        656 => "111011000001",
        657 => "111011000011",
        658 => "111011000100",
        659 => "111011000110",
        660 => "111011001000",
        661 => "111011001001",
        662 => "111011001011",
        663 => "111011001101",
        664 => "111011001110",
        665 => "111011010000",
        666 => "111011010001",
        667 => "111011010011",
        668 => "111011010101",
        669 => "111011010110",
        670 => "111011011000",
        671 => "111011011010",
        672 => "111011011011",
        673 => "111011011101",
        674 => "111011011110",
        675 => "111011100000",
        676 => "111011100010",
        677 => "111011100011",
        678 => "111011100101",
        679 => "111011100110",
        680 => "111011101000",
        681 => "111011101010",
        682 => "111011101011",
        683 => "111011101101",
        684 => "111011101110",
        685 => "111011110000",
        686 => "111011110001",
        687 => "111011110011",
        688 => "111011110101",
        689 => "111011110110",
        690 => "111011111000",
        691 => "111011111001",
        692 => "111011111011",
        693 => "111011111100",
        694 => "111011111110",
        695 => "111011111111",
        696 => "111100000001",
        697 => "111100000010",
        698 => "111100000100",
        699 => "111100000101",
        700 => "111100000111",
        701 => "111100001000",
        702 => "111100001010",
        703 => "111100001011",
        704 => "111100001101",
        705 => "111100001110",
        706 => "111100010000",
        707 => "111100010001",
        708 => "111100010011",
        709 => "111100010100",
        710 => "111100010110",
        711 => "111100010111",
        712 => "111100011000",
        713 => "111100011010",
        714 => "111100011011",
        715 => "111100011101",
        716 => "111100011110",
        717 => "111100100000",
        718 => "111100100001",
        719 => "111100100010",
        720 => "111100100100",
        721 => "111100100101",
        722 => "111100100111",
        723 => "111100101000",
        724 => "111100101001",
        725 => "111100101011",
        726 => "111100101100",
        727 => "111100101110",
        728 => "111100101111",
        729 => "111100110000",
        730 => "111100110010",
        731 => "111100110011",
        732 => "111100110101",
        733 => "111100110110",
        734 => "111100110111",
        735 => "111100111001",
        736 => "111100111010",
        737 => "111100111011",
        738 => "111100111101",
        739 => "111100111110",
        740 => "111100111111",
        741 => "111101000001",
        742 => "111101000010",
        743 => "111101000011",
        744 => "111101000101",
        745 => "111101000110",
        746 => "111101000111",
        747 => "111101001000",
        748 => "111101001010",
        749 => "111101001011",
        750 => "111101001100",
        751 => "111101001110",
        752 => "111101001111",
        753 => "111101010000",
        754 => "111101010001",
        755 => "111101010011",
        756 => "111101010100",
        757 => "111101010101",
        758 => "111101010110",
        759 => "111101011000",
        760 => "111101011001",
        761 => "111101011010",
        762 => "111101011011",
        763 => "111101011101",
        764 => "111101011110",
        765 => "111101011111",
        766 => "111101100000",
        767 => "111101100001",
        768 => "111101100011",
        769 => "111101100100",
        770 => "111101100101",
        771 => "111101100110",
        772 => "111101100111",
        773 => "111101101001",
        774 => "111101101010",
        775 => "111101101011",
        776 => "111101101100",
        777 => "111101101101",
        778 => "111101101110",
        779 => "111101110000",
        780 => "111101110001",
        781 => "111101110010",
        782 => "111101110011",
        783 => "111101110100",
        784 => "111101110101",
        785 => "111101110110",
        786 => "111101111000",
        787 => "111101111001",
        788 => "111101111010",
        789 => "111101111011",
        790 => "111101111100",
        791 => "111101111101",
        792 => "111101111110",
        793 => "111101111111",
        794 => "111110000000",
        795 => "111110000001",
        796 => "111110000011",
        797 => "111110000100",
        798 => "111110000101",
        799 => "111110000110",
        800 => "111110000111",
        801 => "111110001000",
        802 => "111110001001",
        803 => "111110001010",
        804 => "111110001011",
        805 => "111110001100",
        806 => "111110001101",
        807 => "111110001110",
        808 => "111110001111",
        809 => "111110010000",
        810 => "111110010001",
        811 => "111110010010",
        812 => "111110010011",
        813 => "111110010100",
        814 => "111110010101",
        815 => "111110010110",
        816 => "111110010111",
        817 => "111110011000",
        818 => "111110011001",
        819 => "111110011010",
        820 => "111110011011",
        821 => "111110011100",
        822 => "111110011101",
        823 => "111110011110",
        824 => "111110011111",
        825 => "111110100000",
        826 => "111110100001",
        827 => "111110100010",
        828 => "111110100011",
        829 => "111110100100",
        830 => "111110100101",
        831 => "111110100101",
        832 => "111110100110",
        833 => "111110100111",
        834 => "111110101000",
        835 => "111110101001",
        836 => "111110101010",
        837 => "111110101011",
        838 => "111110101100",
        839 => "111110101101",
        840 => "111110101101",
        841 => "111110101110",
        842 => "111110101111",
        843 => "111110110000",
        844 => "111110110001",
        845 => "111110110010",
        846 => "111110110011",
        847 => "111110110011",
        848 => "111110110100",
        849 => "111110110101",
        850 => "111110110110",
        851 => "111110110111",
        852 => "111110111000",
        853 => "111110111000",
        854 => "111110111001",
        855 => "111110111010",
        856 => "111110111011",
        857 => "111110111100",
        858 => "111110111100",
        859 => "111110111101",
        860 => "111110111110",
        861 => "111110111111",
        862 => "111111000000",
        863 => "111111000000",
        864 => "111111000001",
        865 => "111111000010",
        866 => "111111000011",
        867 => "111111000011",
        868 => "111111000100",
        869 => "111111000101",
        870 => "111111000110",
        871 => "111111000110",
        872 => "111111000111",
        873 => "111111001000",
        874 => "111111001001",
        875 => "111111001001",
        876 => "111111001010",
        877 => "111111001011",
        878 => "111111001011",
        879 => "111111001100",
        880 => "111111001101",
        881 => "111111001101",
        882 => "111111001110",
        883 => "111111001111",
        884 => "111111001111",
        885 => "111111010000",
        886 => "111111010001",
        887 => "111111010001",
        888 => "111111010010",
        889 => "111111010011",
        890 => "111111010011",
        891 => "111111010100",
        892 => "111111010101",
        893 => "111111010101",
        894 => "111111010110",
        895 => "111111010111",
        896 => "111111010111",
        897 => "111111011000",
        898 => "111111011000",
        899 => "111111011001",
        900 => "111111011010",
        901 => "111111011010",
        902 => "111111011011",
        903 => "111111011011",
        904 => "111111011100",
        905 => "111111011100",
        906 => "111111011101",
        907 => "111111011110",
        908 => "111111011110",
        909 => "111111011111",
        910 => "111111011111",
        911 => "111111100000",
        912 => "111111100000",
        913 => "111111100001",
        914 => "111111100001",
        915 => "111111100010",
        916 => "111111100010",
        917 => "111111100011",
        918 => "111111100011",
        919 => "111111100100",
        920 => "111111100100",
        921 => "111111100101",
        922 => "111111100101",
        923 => "111111100110",
        924 => "111111100110",
        925 => "111111100111",
        926 => "111111100111",
        927 => "111111101000",
        928 => "111111101000",
        929 => "111111101001",
        930 => "111111101001",
        931 => "111111101010",
        932 => "111111101010",
        933 => "111111101011",
        934 => "111111101011",
        935 => "111111101011",
        936 => "111111101100",
        937 => "111111101100",
        938 => "111111101101",
        939 => "111111101101",
        940 => "111111101110",
        941 => "111111101110",
        942 => "111111101110",
        943 => "111111101111",
        944 => "111111101111",
        945 => "111111101111",
        946 => "111111110000",
        947 => "111111110000",
        948 => "111111110001",
        949 => "111111110001",
        950 => "111111110001",
        951 => "111111110010",
        952 => "111111110010",
        953 => "111111110010",
        954 => "111111110011",
        955 => "111111110011",
        956 => "111111110011",
        957 => "111111110100",
        958 => "111111110100",
        959 => "111111110100",
        960 => "111111110101",
        961 => "111111110101",
        962 => "111111110101",
        963 => "111111110110",
        964 => "111111110110",
        965 => "111111110110",
        966 => "111111110110",
        967 => "111111110111",
        968 => "111111110111",
        969 => "111111110111",
        970 => "111111110111",
        971 => "111111111000",
        972 => "111111111000",
        973 => "111111111000",
        974 => "111111111000",
        975 => "111111111001",
        976 => "111111111001",
        977 => "111111111001",
        978 => "111111111001",
        979 => "111111111010",
        980 => "111111111010",
        981 => "111111111010",
        982 => "111111111010",
        983 => "111111111010",
        984 => "111111111011",
        985 => "111111111011",
        986 => "111111111011",
        987 => "111111111011",
        988 => "111111111011",
        989 => "111111111100",
        990 => "111111111100",
        991 => "111111111100",
        992 => "111111111100",
        993 => "111111111100",
        994 => "111111111100",
        995 => "111111111100",
        996 => "111111111101",
        997 => "111111111101",
        998 => "111111111101",
        999 => "111111111101",
        1000 => "111111111101",
        1001 => "111111111101",
        1002 => "111111111101",
        1003 => "111111111101",
        1004 => "111111111110",
        1005 => "111111111110",
        1006 => "111111111110",
        1007 => "111111111110",
        1008 => "111111111110",
        1009 => "111111111110",
        1010 => "111111111110",
        1011 => "111111111110",
        1012 => "111111111110",
        1013 => "111111111110",
        1014 => "111111111110",
        1015 => "111111111110",
        1016 => "111111111110",
        1017 => "111111111110",
        1018 => "111111111110",
        1019 => "111111111110",
        1020 => "111111111110",
        1021 => "111111111110",
        1022 => "111111111110",
        1023 => "111111111110",
        1024 => "111111111111",
        1025 => "111111111110",
        1026 => "111111111110",
        1027 => "111111111110",
        1028 => "111111111110",
        1029 => "111111111110",
        1030 => "111111111110",
        1031 => "111111111110",
        1032 => "111111111110",
        1033 => "111111111110",
        1034 => "111111111110",
        1035 => "111111111110",
        1036 => "111111111110",
        1037 => "111111111110",
        1038 => "111111111110",
        1039 => "111111111110",
        1040 => "111111111110",
        1041 => "111111111110",
        1042 => "111111111110",
        1043 => "111111111110",
        1044 => "111111111110",
        1045 => "111111111101",
        1046 => "111111111101",
        1047 => "111111111101",
        1048 => "111111111101",
        1049 => "111111111101",
        1050 => "111111111101",
        1051 => "111111111101",
        1052 => "111111111101",
        1053 => "111111111100",
        1054 => "111111111100",
        1055 => "111111111100",
        1056 => "111111111100",
        1057 => "111111111100",
        1058 => "111111111100",
        1059 => "111111111100",
        1060 => "111111111011",
        1061 => "111111111011",
        1062 => "111111111011",
        1063 => "111111111011",
        1064 => "111111111011",
        1065 => "111111111010",
        1066 => "111111111010",
        1067 => "111111111010",
        1068 => "111111111010",
        1069 => "111111111010",
        1070 => "111111111001",
        1071 => "111111111001",
        1072 => "111111111001",
        1073 => "111111111001",
        1074 => "111111111000",
        1075 => "111111111000",
        1076 => "111111111000",
        1077 => "111111111000",
        1078 => "111111110111",
        1079 => "111111110111",
        1080 => "111111110111",
        1081 => "111111110111",
        1082 => "111111110110",
        1083 => "111111110110",
        1084 => "111111110110",
        1085 => "111111110110",
        1086 => "111111110101",
        1087 => "111111110101",
        1088 => "111111110101",
        1089 => "111111110100",
        1090 => "111111110100",
        1091 => "111111110100",
        1092 => "111111110011",
        1093 => "111111110011",
        1094 => "111111110011",
        1095 => "111111110010",
        1096 => "111111110010",
        1097 => "111111110010",
        1098 => "111111110001",
        1099 => "111111110001",
        1100 => "111111110001",
        1101 => "111111110000",
        1102 => "111111110000",
        1103 => "111111101111",
        1104 => "111111101111",
        1105 => "111111101111",
        1106 => "111111101110",
        1107 => "111111101110",
        1108 => "111111101110",
        1109 => "111111101101",
        1110 => "111111101101",
        1111 => "111111101100",
        1112 => "111111101100",
        1113 => "111111101011",
        1114 => "111111101011",
        1115 => "111111101011",
        1116 => "111111101010",
        1117 => "111111101010",
        1118 => "111111101001",
        1119 => "111111101001",
        1120 => "111111101000",
        1121 => "111111101000",
        1122 => "111111100111",
        1123 => "111111100111",
        1124 => "111111100110",
        1125 => "111111100110",
        1126 => "111111100101",
        1127 => "111111100101",
        1128 => "111111100100",
        1129 => "111111100100",
        1130 => "111111100011",
        1131 => "111111100011",
        1132 => "111111100010",
        1133 => "111111100010",
        1134 => "111111100001",
        1135 => "111111100001",
        1136 => "111111100000",
        1137 => "111111100000",
        1138 => "111111011111",
        1139 => "111111011111",
        1140 => "111111011110",
        1141 => "111111011110",
        1142 => "111111011101",
        1143 => "111111011100",
        1144 => "111111011100",
        1145 => "111111011011",
        1146 => "111111011011",
        1147 => "111111011010",
        1148 => "111111011010",
        1149 => "111111011001",
        1150 => "111111011000",
        1151 => "111111011000",
        1152 => "111111010111",
        1153 => "111111010111",
        1154 => "111111010110",
        1155 => "111111010101",
        1156 => "111111010101",
        1157 => "111111010100",
        1158 => "111111010011",
        1159 => "111111010011",
        1160 => "111111010010",
        1161 => "111111010001",
        1162 => "111111010001",
        1163 => "111111010000",
        1164 => "111111001111",
        1165 => "111111001111",
        1166 => "111111001110",
        1167 => "111111001101",
        1168 => "111111001101",
        1169 => "111111001100",
        1170 => "111111001011",
        1171 => "111111001011",
        1172 => "111111001010",
        1173 => "111111001001",
        1174 => "111111001001",
        1175 => "111111001000",
        1176 => "111111000111",
        1177 => "111111000110",
        1178 => "111111000110",
        1179 => "111111000101",
        1180 => "111111000100",
        1181 => "111111000011",
        1182 => "111111000011",
        1183 => "111111000010",
        1184 => "111111000001",
        1185 => "111111000000",
        1186 => "111111000000",
        1187 => "111110111111",
        1188 => "111110111110",
        1189 => "111110111101",
        1190 => "111110111100",
        1191 => "111110111100",
        1192 => "111110111011",
        1193 => "111110111010",
        1194 => "111110111001",
        1195 => "111110111000",
        1196 => "111110111000",
        1197 => "111110110111",
        1198 => "111110110110",
        1199 => "111110110101",
        1200 => "111110110100",
        1201 => "111110110011",
        1202 => "111110110011",
        1203 => "111110110010",
        1204 => "111110110001",
        1205 => "111110110000",
        1206 => "111110101111",
        1207 => "111110101110",
        1208 => "111110101101",
        1209 => "111110101101",
        1210 => "111110101100",
        1211 => "111110101011",
        1212 => "111110101010",
        1213 => "111110101001",
        1214 => "111110101000",
        1215 => "111110100111",
        1216 => "111110100110",
        1217 => "111110100101",
        1218 => "111110100101",
        1219 => "111110100100",
        1220 => "111110100011",
        1221 => "111110100010",
        1222 => "111110100001",
        1223 => "111110100000",
        1224 => "111110011111",
        1225 => "111110011110",
        1226 => "111110011101",
        1227 => "111110011100",
        1228 => "111110011011",
        1229 => "111110011010",
        1230 => "111110011001",
        1231 => "111110011000",
        1232 => "111110010111",
        1233 => "111110010110",
        1234 => "111110010101",
        1235 => "111110010100",
        1236 => "111110010011",
        1237 => "111110010010",
        1238 => "111110010001",
        1239 => "111110010000",
        1240 => "111110001111",
        1241 => "111110001110",
        1242 => "111110001101",
        1243 => "111110001100",
        1244 => "111110001011",
        1245 => "111110001010",
        1246 => "111110001001",
        1247 => "111110001000",
        1248 => "111110000111",
        1249 => "111110000110",
        1250 => "111110000101",
        1251 => "111110000100",
        1252 => "111110000011",
        1253 => "111110000001",
        1254 => "111110000000",
        1255 => "111101111111",
        1256 => "111101111110",
        1257 => "111101111101",
        1258 => "111101111100",
        1259 => "111101111011",
        1260 => "111101111010",
        1261 => "111101111001",
        1262 => "111101111000",
        1263 => "111101110110",
        1264 => "111101110101",
        1265 => "111101110100",
        1266 => "111101110011",
        1267 => "111101110010",
        1268 => "111101110001",
        1269 => "111101110000",
        1270 => "111101101110",
        1271 => "111101101101",
        1272 => "111101101100",
        1273 => "111101101011",
        1274 => "111101101010",
        1275 => "111101101001",
        1276 => "111101100111",
        1277 => "111101100110",
        1278 => "111101100101",
        1279 => "111101100100",
        1280 => "111101100011",
        1281 => "111101100001",
        1282 => "111101100000",
        1283 => "111101011111",
        1284 => "111101011110",
        1285 => "111101011101",
        1286 => "111101011011",
        1287 => "111101011010",
        1288 => "111101011001",
        1289 => "111101011000",
        1290 => "111101010110",
        1291 => "111101010101",
        1292 => "111101010100",
        1293 => "111101010011",
        1294 => "111101010001",
        1295 => "111101010000",
        1296 => "111101001111",
        1297 => "111101001110",
        1298 => "111101001100",
        1299 => "111101001011",
        1300 => "111101001010",
        1301 => "111101001000",
        1302 => "111101000111",
        1303 => "111101000110",
        1304 => "111101000101",
        1305 => "111101000011",
        1306 => "111101000010",
        1307 => "111101000001",
        1308 => "111100111111",
        1309 => "111100111110",
        1310 => "111100111101",
        1311 => "111100111011",
        1312 => "111100111010",
        1313 => "111100111001",
        1314 => "111100110111",
        1315 => "111100110110",
        1316 => "111100110101",
        1317 => "111100110011",
        1318 => "111100110010",
        1319 => "111100110000",
        1320 => "111100101111",
        1321 => "111100101110",
        1322 => "111100101100",
        1323 => "111100101011",
        1324 => "111100101001",
        1325 => "111100101000",
        1326 => "111100100111",
        1327 => "111100100101",
        1328 => "111100100100",
        1329 => "111100100010",
        1330 => "111100100001",
        1331 => "111100100000",
        1332 => "111100011110",
        1333 => "111100011101",
        1334 => "111100011011",
        1335 => "111100011010",
        1336 => "111100011000",
        1337 => "111100010111",
        1338 => "111100010110",
        1339 => "111100010100",
        1340 => "111100010011",
        1341 => "111100010001",
        1342 => "111100010000",
        1343 => "111100001110",
        1344 => "111100001101",
        1345 => "111100001011",
        1346 => "111100001010",
        1347 => "111100001000",
        1348 => "111100000111",
        1349 => "111100000101",
        1350 => "111100000100",
        1351 => "111100000010",
        1352 => "111100000001",
        1353 => "111011111111",
        1354 => "111011111110",
        1355 => "111011111100",
        1356 => "111011111011",
        1357 => "111011111001",
        1358 => "111011111000",
        1359 => "111011110110",
        1360 => "111011110101",
        1361 => "111011110011",
        1362 => "111011110001",
        1363 => "111011110000",
        1364 => "111011101110",
        1365 => "111011101101",
        1366 => "111011101011",
        1367 => "111011101010",
        1368 => "111011101000",
        1369 => "111011100110",
        1370 => "111011100101",
        1371 => "111011100011",
        1372 => "111011100010",
        1373 => "111011100000",
        1374 => "111011011110",
        1375 => "111011011101",
        1376 => "111011011011",
        1377 => "111011011010",
        1378 => "111011011000",
        1379 => "111011010110",
        1380 => "111011010101",
        1381 => "111011010011",
        1382 => "111011010001",
        1383 => "111011010000",
        1384 => "111011001110",
        1385 => "111011001101",
        1386 => "111011001011",
        1387 => "111011001001",
        1388 => "111011001000",
        1389 => "111011000110",
        1390 => "111011000100",
        1391 => "111011000011",
        1392 => "111011000001",
        1393 => "111010111111",
        1394 => "111010111101",
        1395 => "111010111100",
        1396 => "111010111010",
        1397 => "111010111000",
        1398 => "111010110111",
        1399 => "111010110101",
        1400 => "111010110011",
        1401 => "111010110010",
        1402 => "111010110000",
        1403 => "111010101110",
        1404 => "111010101100",
        1405 => "111010101011",
        1406 => "111010101001",
        1407 => "111010100111",
        1408 => "111010100101",
        1409 => "111010100100",
        1410 => "111010100010",
        1411 => "111010100000",
        1412 => "111010011110",
        1413 => "111010011101",
        1414 => "111010011011",
        1415 => "111010011001",
        1416 => "111010010111",
        1417 => "111010010110",
        1418 => "111010010100",
        1419 => "111010010010",
        1420 => "111010010000",
        1421 => "111010001110",
        1422 => "111010001101",
        1423 => "111010001011",
        1424 => "111010001001",
        1425 => "111010000111",
        1426 => "111010000101",
        1427 => "111010000100",
        1428 => "111010000010",
        1429 => "111010000000",
        1430 => "111001111110",
        1431 => "111001111100",
        1432 => "111001111010",
        1433 => "111001111001",
        1434 => "111001110111",
        1435 => "111001110101",
        1436 => "111001110011",
        1437 => "111001110001",
        1438 => "111001101111",
        1439 => "111001101101",
        1440 => "111001101100",
        1441 => "111001101010",
        1442 => "111001101000",
        1443 => "111001100110",
        1444 => "111001100100",
        1445 => "111001100010",
        1446 => "111001100000",
        1447 => "111001011110",
        1448 => "111001011100",
        1449 => "111001011011",
        1450 => "111001011001",
        1451 => "111001010111",
        1452 => "111001010101",
        1453 => "111001010011",
        1454 => "111001010001",
        1455 => "111001001111",
        1456 => "111001001101",
        1457 => "111001001011",
        1458 => "111001001001",
        1459 => "111001000111",
        1460 => "111001000101",
        1461 => "111001000011",
        1462 => "111001000001",
        1463 => "111001000000",
        1464 => "111000111110",
        1465 => "111000111100",
        1466 => "111000111010",
        1467 => "111000111000",
        1468 => "111000110110",
        1469 => "111000110100",
        1470 => "111000110010",
        1471 => "111000110000",
        1472 => "111000101110",
        1473 => "111000101100",
        1474 => "111000101010",
        1475 => "111000101000",
        1476 => "111000100110",
        1477 => "111000100100",
        1478 => "111000100010",
        1479 => "111000100000",
        1480 => "111000011110",
        1481 => "111000011100",
        1482 => "111000011010",
        1483 => "111000011000",
        1484 => "111000010110",
        1485 => "111000010100",
        1486 => "111000010001",
        1487 => "111000001111",
        1488 => "111000001101",
        1489 => "111000001011",
        1490 => "111000001001",
        1491 => "111000000111",
        1492 => "111000000101",
        1493 => "111000000011",
        1494 => "111000000001",
        1495 => "110111111111",
        1496 => "110111111101",
        1497 => "110111111011",
        1498 => "110111111001",
        1499 => "110111110111",
        1500 => "110111110101",
        1501 => "110111110010",
        1502 => "110111110000",
        1503 => "110111101110",
        1504 => "110111101100",
        1505 => "110111101010",
        1506 => "110111101000",
        1507 => "110111100110",
        1508 => "110111100100",
        1509 => "110111100010",
        1510 => "110111011111",
        1511 => "110111011101",
        1512 => "110111011011",
        1513 => "110111011001",
        1514 => "110111010111",
        1515 => "110111010101",
        1516 => "110111010011",
        1517 => "110111010000",
        1518 => "110111001110",
        1519 => "110111001100",
        1520 => "110111001010",
        1521 => "110111001000",
        1522 => "110111000110",
        1523 => "110111000011",
        1524 => "110111000001",
        1525 => "110110111111",
        1526 => "110110111101",
        1527 => "110110111011",
        1528 => "110110111000",
        1529 => "110110110110",
        1530 => "110110110100",
        1531 => "110110110010",
        1532 => "110110110000",
        1533 => "110110101101",
        1534 => "110110101011",
        1535 => "110110101001",
        1536 => "110110100111",
        1537 => "110110100101",
        1538 => "110110100010",
        1539 => "110110100000",
        1540 => "110110011110",
        1541 => "110110011100",
        1542 => "110110011001",
        1543 => "110110010111",
        1544 => "110110010101",
        1545 => "110110010011",
        1546 => "110110010000",
        1547 => "110110001110",
        1548 => "110110001100",
        1549 => "110110001010",
        1550 => "110110000111",
        1551 => "110110000101",
        1552 => "110110000011",
        1553 => "110110000001",
        1554 => "110101111110",
        1555 => "110101111100",
        1556 => "110101111010",
        1557 => "110101110111",
        1558 => "110101110101",
        1559 => "110101110011",
        1560 => "110101110001",
        1561 => "110101101110",
        1562 => "110101101100",
        1563 => "110101101010",
        1564 => "110101100111",
        1565 => "110101100101",
        1566 => "110101100011",
        1567 => "110101100000",
        1568 => "110101011110",
        1569 => "110101011100",
        1570 => "110101011001",
        1571 => "110101010111",
        1572 => "110101010101",
        1573 => "110101010010",
        1574 => "110101010000",
        1575 => "110101001110",
        1576 => "110101001011",
        1577 => "110101001001",
        1578 => "110101000111",
        1579 => "110101000100",
        1580 => "110101000010",
        1581 => "110100111111",
        1582 => "110100111101",
        1583 => "110100111011",
        1584 => "110100111000",
        1585 => "110100110110",
        1586 => "110100110100",
        1587 => "110100110001",
        1588 => "110100101111",
        1589 => "110100101100",
        1590 => "110100101010",
        1591 => "110100101000",
        1592 => "110100100101",
        1593 => "110100100011",
        1594 => "110100100000",
        1595 => "110100011110",
        1596 => "110100011100",
        1597 => "110100011001",
        1598 => "110100010111",
        1599 => "110100010100",
        1600 => "110100010010",
        1601 => "110100001111",
        1602 => "110100001101",
        1603 => "110100001011",
        1604 => "110100001000",
        1605 => "110100000110",
        1606 => "110100000011",
        1607 => "110100000001",
        1608 => "110011111110",
        1609 => "110011111100",
        1610 => "110011111001",
        1611 => "110011110111",
        1612 => "110011110101",
        1613 => "110011110010",
        1614 => "110011110000",
        1615 => "110011101101",
        1616 => "110011101011",
        1617 => "110011101000",
        1618 => "110011100110",
        1619 => "110011100011",
        1620 => "110011100001",
        1621 => "110011011110",
        1622 => "110011011100",
        1623 => "110011011001",
        1624 => "110011010111",
        1625 => "110011010100",
        1626 => "110011010010",
        1627 => "110011001111",
        1628 => "110011001101",
        1629 => "110011001010",
        1630 => "110011001000",
        1631 => "110011000101",
        1632 => "110011000011",
        1633 => "110011000000",
        1634 => "110010111110",
        1635 => "110010111011",
        1636 => "110010111001",
        1637 => "110010110110",
        1638 => "110010110100",
        1639 => "110010110001",
        1640 => "110010101110",
        1641 => "110010101100",
        1642 => "110010101001",
        1643 => "110010100111",
        1644 => "110010100100",
        1645 => "110010100010",
        1646 => "110010011111",
        1647 => "110010011101",
        1648 => "110010011010",
        1649 => "110010010111",
        1650 => "110010010101",
        1651 => "110010010010",
        1652 => "110010010000",
        1653 => "110010001101",
        1654 => "110010001011",
        1655 => "110010001000",
        1656 => "110010000101",
        1657 => "110010000011",
        1658 => "110010000000",
        1659 => "110001111110",
        1660 => "110001111011",
        1661 => "110001111000",
        1662 => "110001110110",
        1663 => "110001110011",
        1664 => "110001110001",
        1665 => "110001101110",
        1666 => "110001101011",
        1667 => "110001101001",
        1668 => "110001100110",
        1669 => "110001100011",
        1670 => "110001100001",
        1671 => "110001011110",
        1672 => "110001011100",
        1673 => "110001011001",
        1674 => "110001010110",
        1675 => "110001010100",
        1676 => "110001010001",
        1677 => "110001001110",
        1678 => "110001001100",
        1679 => "110001001001",
        1680 => "110001000110",
        1681 => "110001000100",
        1682 => "110001000001",
        1683 => "110000111110",
        1684 => "110000111100",
        1685 => "110000111001",
        1686 => "110000110110",
        1687 => "110000110100",
        1688 => "110000110001",
        1689 => "110000101110",
        1690 => "110000101100",
        1691 => "110000101001",
        1692 => "110000100110",
        1693 => "110000100100",
        1694 => "110000100001",
        1695 => "110000011110",
        1696 => "110000011100",
        1697 => "110000011001",
        1698 => "110000010110",
        1699 => "110000010100",
        1700 => "110000010001",
        1701 => "110000001110",
        1702 => "110000001011",
        1703 => "110000001001",
        1704 => "110000000110",
        1705 => "110000000011",
        1706 => "110000000001",
        1707 => "101111111110",
        1708 => "101111111011",
        1709 => "101111111000",
        1710 => "101111110110",
        1711 => "101111110011",
        1712 => "101111110000",
        1713 => "101111101101",
        1714 => "101111101011",
        1715 => "101111101000",
        1716 => "101111100101",
        1717 => "101111100011",
        1718 => "101111100000",
        1719 => "101111011101",
        1720 => "101111011010",
        1721 => "101111011000",
        1722 => "101111010101",
        1723 => "101111010010",
        1724 => "101111001111",
        1725 => "101111001100",
        1726 => "101111001010",
        1727 => "101111000111",
        1728 => "101111000100",
        1729 => "101111000001",
        1730 => "101110111111",
        1731 => "101110111100",
        1732 => "101110111001",
        1733 => "101110110110",
        1734 => "101110110100",
        1735 => "101110110001",
        1736 => "101110101110",
        1737 => "101110101011",
        1738 => "101110101000",
        1739 => "101110100110",
        1740 => "101110100011",
        1741 => "101110100000",
        1742 => "101110011101",
        1743 => "101110011010",
        1744 => "101110011000",
        1745 => "101110010101",
        1746 => "101110010010",
        1747 => "101110001111",
        1748 => "101110001100",
        1749 => "101110001010",
        1750 => "101110000111",
        1751 => "101110000100",
        1752 => "101110000001",
        1753 => "101101111110",
        1754 => "101101111011",
        1755 => "101101111001",
        1756 => "101101110110",
        1757 => "101101110011",
        1758 => "101101110000",
        1759 => "101101101101",
        1760 => "101101101010",
        1761 => "101101101000",
        1762 => "101101100101",
        1763 => "101101100010",
        1764 => "101101011111",
        1765 => "101101011100",
        1766 => "101101011001",
        1767 => "101101010110",
        1768 => "101101010100",
        1769 => "101101010001",
        1770 => "101101001110",
        1771 => "101101001011",
        1772 => "101101001000",
        1773 => "101101000101",
        1774 => "101101000010",
        1775 => "101101000000",
        1776 => "101100111101",
        1777 => "101100111010",
        1778 => "101100110111",
        1779 => "101100110100",
        1780 => "101100110001",
        1781 => "101100101110",
        1782 => "101100101011",
        1783 => "101100101001",
        1784 => "101100100110",
        1785 => "101100100011",
        1786 => "101100100000",
        1787 => "101100011101",
        1788 => "101100011010",
        1789 => "101100010111",
        1790 => "101100010100",
        1791 => "101100010001",
        1792 => "101100001111",
        1793 => "101100001100",
        1794 => "101100001001",
        1795 => "101100000110",
        1796 => "101100000011",
        1797 => "101100000000",
        1798 => "101011111101",
        1799 => "101011111010",
        1800 => "101011110111",
        1801 => "101011110100",
        1802 => "101011110001",
        1803 => "101011101111",
        1804 => "101011101100",
        1805 => "101011101001",
        1806 => "101011100110",
        1807 => "101011100011",
        1808 => "101011100000",
        1809 => "101011011101",
        1810 => "101011011010",
        1811 => "101011010111",
        1812 => "101011010100",
        1813 => "101011010001",
        1814 => "101011001110",
        1815 => "101011001011",
        1816 => "101011001000",
        1817 => "101011000101",
        1818 => "101011000010",
        1819 => "101011000000",
        1820 => "101010111101",
        1821 => "101010111010",
        1822 => "101010110111",
        1823 => "101010110100",
        1824 => "101010110001",
        1825 => "101010101110",
        1826 => "101010101011",
        1827 => "101010101000",
        1828 => "101010100101",
        1829 => "101010100010",
        1830 => "101010011111",
        1831 => "101010011100",
        1832 => "101010011001",
        1833 => "101010010110",
        1834 => "101010010011",
        1835 => "101010010000",
        1836 => "101010001101",
        1837 => "101010001010",
        1838 => "101010000111",
        1839 => "101010000100",
        1840 => "101010000001",
        1841 => "101001111110",
        1842 => "101001111011",
        1843 => "101001111000",
        1844 => "101001110101",
        1845 => "101001110010",
        1846 => "101001101111",
        1847 => "101001101100",
        1848 => "101001101001",
        1849 => "101001100110",
        1850 => "101001100011",
        1851 => "101001100000",
        1852 => "101001011101",
        1853 => "101001011010",
        1854 => "101001010111",
        1855 => "101001010100",
        1856 => "101001010001",
        1857 => "101001001110",
        1858 => "101001001011",
        1859 => "101001001000",
        1860 => "101001000101",
        1861 => "101001000010",
        1862 => "101000111111",
        1863 => "101000111100",
        1864 => "101000111001",
        1865 => "101000110110",
        1866 => "101000110011",
        1867 => "101000110000",
        1868 => "101000101101",
        1869 => "101000101010",
        1870 => "101000100111",
        1871 => "101000100100",
        1872 => "101000100001",
        1873 => "101000011110",
        1874 => "101000011011",
        1875 => "101000011000",
        1876 => "101000010101",
        1877 => "101000010010",
        1878 => "101000001111",
        1879 => "101000001100",
        1880 => "101000001001",
        1881 => "101000000110",
        1882 => "101000000011",
        1883 => "101000000000",
        1884 => "100111111101",
        1885 => "100111111010",
        1886 => "100111110111",
        1887 => "100111110100",
        1888 => "100111110001",
        1889 => "100111101101",
        1890 => "100111101010",
        1891 => "100111100111",
        1892 => "100111100100",
        1893 => "100111100001",
        1894 => "100111011110",
        1895 => "100111011011",
        1896 => "100111011000",
        1897 => "100111010101",
        1898 => "100111010010",
        1899 => "100111001111",
        1900 => "100111001100",
        1901 => "100111001001",
        1902 => "100111000110",
        1903 => "100111000011",
        1904 => "100111000000",
        1905 => "100110111101",
        1906 => "100110111001",
        1907 => "100110110110",
        1908 => "100110110011",
        1909 => "100110110000",
        1910 => "100110101101",
        1911 => "100110101010",
        1912 => "100110100111",
        1913 => "100110100100",
        1914 => "100110100001",
        1915 => "100110011110",
        1916 => "100110011011",
        1917 => "100110011000",
        1918 => "100110010101",
        1919 => "100110010010",
        1920 => "100110001110",
        1921 => "100110001011",
        1922 => "100110001000",
        1923 => "100110000101",
        1924 => "100110000010",
        1925 => "100101111111",
        1926 => "100101111100",
        1927 => "100101111001",
        1928 => "100101110110",
        1929 => "100101110011",
        1930 => "100101110000",
        1931 => "100101101101",
        1932 => "100101101001",
        1933 => "100101100110",
        1934 => "100101100011",
        1935 => "100101100000",
        1936 => "100101011101",
        1937 => "100101011010",
        1938 => "100101010111",
        1939 => "100101010100",
        1940 => "100101010001",
        1941 => "100101001110",
        1942 => "100101001010",
        1943 => "100101000111",
        1944 => "100101000100",
        1945 => "100101000001",
        1946 => "100100111110",
        1947 => "100100111011",
        1948 => "100100111000",
        1949 => "100100110101",
        1950 => "100100110010",
        1951 => "100100101111",
        1952 => "100100101011",
        1953 => "100100101000",
        1954 => "100100100101",
        1955 => "100100100010",
        1956 => "100100011111",
        1957 => "100100011100",
        1958 => "100100011001",
        1959 => "100100010110",
        1960 => "100100010011",
        1961 => "100100001111",
        1962 => "100100001100",
        1963 => "100100001001",
        1964 => "100100000110",
        1965 => "100100000011",
        1966 => "100100000000",
        1967 => "100011111101",
        1968 => "100011111010",
        1969 => "100011110111",
        1970 => "100011110011",
        1971 => "100011110000",
        1972 => "100011101101",
        1973 => "100011101010",
        1974 => "100011100111",
        1975 => "100011100100",
        1976 => "100011100001",
        1977 => "100011011110",
        1978 => "100011011010",
        1979 => "100011010111",
        1980 => "100011010100",
        1981 => "100011010001",
        1982 => "100011001110",
        1983 => "100011001011",
        1984 => "100011001000",
        1985 => "100011000101",
        1986 => "100011000001",
        1987 => "100010111110",
        1988 => "100010111011",
        1989 => "100010111000",
        1990 => "100010110101",
        1991 => "100010110010",
        1992 => "100010101111",
        1993 => "100010101100",
        1994 => "100010101000",
        1995 => "100010100101",
        1996 => "100010100010",
        1997 => "100010011111",
        1998 => "100010011100",
        1999 => "100010011001",
        2000 => "100010010110",
        2001 => "100010010010",
        2002 => "100010001111",
        2003 => "100010001100",
        2004 => "100010001001",
        2005 => "100010000110",
        2006 => "100010000011",
        2007 => "100010000000",
        2008 => "100001111101",
        2009 => "100001111001",
        2010 => "100001110110",
        2011 => "100001110011",
        2012 => "100001110000",
        2013 => "100001101101",
        2014 => "100001101010",
        2015 => "100001100111",
        2016 => "100001100011",
        2017 => "100001100000",
        2018 => "100001011101",
        2019 => "100001011010",
        2020 => "100001010111",
        2021 => "100001010100",
        2022 => "100001010001",
        2023 => "100001001110",
        2024 => "100001001010",
        2025 => "100001000111",
        2026 => "100001000100",
        2027 => "100001000001",
        2028 => "100000111110",
        2029 => "100000111011",
        2030 => "100000111000",
        2031 => "100000110100",
        2032 => "100000110001",
        2033 => "100000101110",
        2034 => "100000101011",
        2035 => "100000101000",
        2036 => "100000100101",
        2037 => "100000100010",
        2038 => "100000011110",
        2039 => "100000011011",
        2040 => "100000011000",
        2041 => "100000010101",
        2042 => "100000010010",
        2043 => "100000001111",
        2044 => "100000001100",
        2045 => "100000001000",
        2046 => "100000000101",
        2047 => "100000000010",
        2048 => "011111111111",
        2049 => "011111111100",
        2050 => "011111111001",
        2051 => "011111110110",
        2052 => "011111110010",
        2053 => "011111101111",
        2054 => "011111101100",
        2055 => "011111101001",
        2056 => "011111100110",
        2057 => "011111100011",
        2058 => "011111100000",
        2059 => "011111011100",
        2060 => "011111011001",
        2061 => "011111010110",
        2062 => "011111010011",
        2063 => "011111010000",
        2064 => "011111001101",
        2065 => "011111001010",
        2066 => "011111000110",
        2067 => "011111000011",
        2068 => "011111000000",
        2069 => "011110111101",
        2070 => "011110111010",
        2071 => "011110110111",
        2072 => "011110110100",
        2073 => "011110110000",
        2074 => "011110101101",
        2075 => "011110101010",
        2076 => "011110100111",
        2077 => "011110100100",
        2078 => "011110100001",
        2079 => "011110011110",
        2080 => "011110011011",
        2081 => "011110010111",
        2082 => "011110010100",
        2083 => "011110010001",
        2084 => "011110001110",
        2085 => "011110001011",
        2086 => "011110001000",
        2087 => "011110000101",
        2088 => "011110000001",
        2089 => "011101111110",
        2090 => "011101111011",
        2091 => "011101111000",
        2092 => "011101110101",
        2093 => "011101110010",
        2094 => "011101101111",
        2095 => "011101101100",
        2096 => "011101101000",
        2097 => "011101100101",
        2098 => "011101100010",
        2099 => "011101011111",
        2100 => "011101011100",
        2101 => "011101011001",
        2102 => "011101010110",
        2103 => "011101010010",
        2104 => "011101001111",
        2105 => "011101001100",
        2106 => "011101001001",
        2107 => "011101000110",
        2108 => "011101000011",
        2109 => "011101000000",
        2110 => "011100111101",
        2111 => "011100111001",
        2112 => "011100110110",
        2113 => "011100110011",
        2114 => "011100110000",
        2115 => "011100101101",
        2116 => "011100101010",
        2117 => "011100100111",
        2118 => "011100100100",
        2119 => "011100100000",
        2120 => "011100011101",
        2121 => "011100011010",
        2122 => "011100010111",
        2123 => "011100010100",
        2124 => "011100010001",
        2125 => "011100001110",
        2126 => "011100001011",
        2127 => "011100000111",
        2128 => "011100000100",
        2129 => "011100000001",
        2130 => "011011111110",
        2131 => "011011111011",
        2132 => "011011111000",
        2133 => "011011110101",
        2134 => "011011110010",
        2135 => "011011101111",
        2136 => "011011101011",
        2137 => "011011101000",
        2138 => "011011100101",
        2139 => "011011100010",
        2140 => "011011011111",
        2141 => "011011011100",
        2142 => "011011011001",
        2143 => "011011010110",
        2144 => "011011010011",
        2145 => "011011001111",
        2146 => "011011001100",
        2147 => "011011001001",
        2148 => "011011000110",
        2149 => "011011000011",
        2150 => "011011000000",
        2151 => "011010111101",
        2152 => "011010111010",
        2153 => "011010110111",
        2154 => "011010110100",
        2155 => "011010110000",
        2156 => "011010101101",
        2157 => "011010101010",
        2158 => "011010100111",
        2159 => "011010100100",
        2160 => "011010100001",
        2161 => "011010011110",
        2162 => "011010011011",
        2163 => "011010011000",
        2164 => "011010010101",
        2165 => "011010010001",
        2166 => "011010001110",
        2167 => "011010001011",
        2168 => "011010001000",
        2169 => "011010000101",
        2170 => "011010000010",
        2171 => "011001111111",
        2172 => "011001111100",
        2173 => "011001111001",
        2174 => "011001110110",
        2175 => "011001110011",
        2176 => "011001110000",
        2177 => "011001101100",
        2178 => "011001101001",
        2179 => "011001100110",
        2180 => "011001100011",
        2181 => "011001100000",
        2182 => "011001011101",
        2183 => "011001011010",
        2184 => "011001010111",
        2185 => "011001010100",
        2186 => "011001010001",
        2187 => "011001001110",
        2188 => "011001001011",
        2189 => "011001001000",
        2190 => "011001000101",
        2191 => "011001000001",
        2192 => "011000111110",
        2193 => "011000111011",
        2194 => "011000111000",
        2195 => "011000110101",
        2196 => "011000110010",
        2197 => "011000101111",
        2198 => "011000101100",
        2199 => "011000101001",
        2200 => "011000100110",
        2201 => "011000100011",
        2202 => "011000100000",
        2203 => "011000011101",
        2204 => "011000011010",
        2205 => "011000010111",
        2206 => "011000010100",
        2207 => "011000010001",
        2208 => "011000001101",
        2209 => "011000001010",
        2210 => "011000000111",
        2211 => "011000000100",
        2212 => "011000000001",
        2213 => "010111111110",
        2214 => "010111111011",
        2215 => "010111111000",
        2216 => "010111110101",
        2217 => "010111110010",
        2218 => "010111101111",
        2219 => "010111101100",
        2220 => "010111101001",
        2221 => "010111100110",
        2222 => "010111100011",
        2223 => "010111100000",
        2224 => "010111011101",
        2225 => "010111011010",
        2226 => "010111010111",
        2227 => "010111010100",
        2228 => "010111010001",
        2229 => "010111001110",
        2230 => "010111001011",
        2231 => "010111001000",
        2232 => "010111000101",
        2233 => "010111000010",
        2234 => "010110111111",
        2235 => "010110111100",
        2236 => "010110111001",
        2237 => "010110110110",
        2238 => "010110110011",
        2239 => "010110110000",
        2240 => "010110101101",
        2241 => "010110101010",
        2242 => "010110100111",
        2243 => "010110100100",
        2244 => "010110100001",
        2245 => "010110011110",
        2246 => "010110011011",
        2247 => "010110011000",
        2248 => "010110010101",
        2249 => "010110010010",
        2250 => "010110001111",
        2251 => "010110001100",
        2252 => "010110001001",
        2253 => "010110000110",
        2254 => "010110000011",
        2255 => "010110000000",
        2256 => "010101111101",
        2257 => "010101111010",
        2258 => "010101110111",
        2259 => "010101110100",
        2260 => "010101110001",
        2261 => "010101101110",
        2262 => "010101101011",
        2263 => "010101101000",
        2264 => "010101100101",
        2265 => "010101100010",
        2266 => "010101011111",
        2267 => "010101011100",
        2268 => "010101011001",
        2269 => "010101010110",
        2270 => "010101010011",
        2271 => "010101010000",
        2272 => "010101001101",
        2273 => "010101001010",
        2274 => "010101000111",
        2275 => "010101000100",
        2276 => "010101000001",
        2277 => "010100111110",
        2278 => "010100111100",
        2279 => "010100111001",
        2280 => "010100110110",
        2281 => "010100110011",
        2282 => "010100110000",
        2283 => "010100101101",
        2284 => "010100101010",
        2285 => "010100100111",
        2286 => "010100100100",
        2287 => "010100100001",
        2288 => "010100011110",
        2289 => "010100011011",
        2290 => "010100011000",
        2291 => "010100010101",
        2292 => "010100010010",
        2293 => "010100001111",
        2294 => "010100001101",
        2295 => "010100001010",
        2296 => "010100000111",
        2297 => "010100000100",
        2298 => "010100000001",
        2299 => "010011111110",
        2300 => "010011111011",
        2301 => "010011111000",
        2302 => "010011110101",
        2303 => "010011110010",
        2304 => "010011101111",
        2305 => "010011101101",
        2306 => "010011101010",
        2307 => "010011100111",
        2308 => "010011100100",
        2309 => "010011100001",
        2310 => "010011011110",
        2311 => "010011011011",
        2312 => "010011011000",
        2313 => "010011010101",
        2314 => "010011010011",
        2315 => "010011010000",
        2316 => "010011001101",
        2317 => "010011001010",
        2318 => "010011000111",
        2319 => "010011000100",
        2320 => "010011000001",
        2321 => "010010111110",
        2322 => "010010111100",
        2323 => "010010111001",
        2324 => "010010110110",
        2325 => "010010110011",
        2326 => "010010110000",
        2327 => "010010101101",
        2328 => "010010101010",
        2329 => "010010101000",
        2330 => "010010100101",
        2331 => "010010100010",
        2332 => "010010011111",
        2333 => "010010011100",
        2334 => "010010011001",
        2335 => "010010010110",
        2336 => "010010010100",
        2337 => "010010010001",
        2338 => "010010001110",
        2339 => "010010001011",
        2340 => "010010001000",
        2341 => "010010000101",
        2342 => "010010000011",
        2343 => "010010000000",
        2344 => "010001111101",
        2345 => "010001111010",
        2346 => "010001110111",
        2347 => "010001110100",
        2348 => "010001110010",
        2349 => "010001101111",
        2350 => "010001101100",
        2351 => "010001101001",
        2352 => "010001100110",
        2353 => "010001100100",
        2354 => "010001100001",
        2355 => "010001011110",
        2356 => "010001011011",
        2357 => "010001011000",
        2358 => "010001010110",
        2359 => "010001010011",
        2360 => "010001010000",
        2361 => "010001001101",
        2362 => "010001001010",
        2363 => "010001001000",
        2364 => "010001000101",
        2365 => "010001000010",
        2366 => "010000111111",
        2367 => "010000111101",
        2368 => "010000111010",
        2369 => "010000110111",
        2370 => "010000110100",
        2371 => "010000110010",
        2372 => "010000101111",
        2373 => "010000101100",
        2374 => "010000101001",
        2375 => "010000100110",
        2376 => "010000100100",
        2377 => "010000100001",
        2378 => "010000011110",
        2379 => "010000011011",
        2380 => "010000011001",
        2381 => "010000010110",
        2382 => "010000010011",
        2383 => "010000010001",
        2384 => "010000001110",
        2385 => "010000001011",
        2386 => "010000001000",
        2387 => "010000000110",
        2388 => "010000000011",
        2389 => "010000000000",
        2390 => "001111111101",
        2391 => "001111111011",
        2392 => "001111111000",
        2393 => "001111110101",
        2394 => "001111110011",
        2395 => "001111110000",
        2396 => "001111101101",
        2397 => "001111101010",
        2398 => "001111101000",
        2399 => "001111100101",
        2400 => "001111100010",
        2401 => "001111100000",
        2402 => "001111011101",
        2403 => "001111011010",
        2404 => "001111011000",
        2405 => "001111010101",
        2406 => "001111010010",
        2407 => "001111010000",
        2408 => "001111001101",
        2409 => "001111001010",
        2410 => "001111001000",
        2411 => "001111000101",
        2412 => "001111000010",
        2413 => "001111000000",
        2414 => "001110111101",
        2415 => "001110111010",
        2416 => "001110111000",
        2417 => "001110110101",
        2418 => "001110110010",
        2419 => "001110110000",
        2420 => "001110101101",
        2421 => "001110101010",
        2422 => "001110101000",
        2423 => "001110100101",
        2424 => "001110100010",
        2425 => "001110100000",
        2426 => "001110011101",
        2427 => "001110011011",
        2428 => "001110011000",
        2429 => "001110010101",
        2430 => "001110010011",
        2431 => "001110010000",
        2432 => "001110001101",
        2433 => "001110001011",
        2434 => "001110001000",
        2435 => "001110000110",
        2436 => "001110000011",
        2437 => "001110000000",
        2438 => "001101111110",
        2439 => "001101111011",
        2440 => "001101111001",
        2441 => "001101110110",
        2442 => "001101110011",
        2443 => "001101110001",
        2444 => "001101101110",
        2445 => "001101101100",
        2446 => "001101101001",
        2447 => "001101100111",
        2448 => "001101100100",
        2449 => "001101100001",
        2450 => "001101011111",
        2451 => "001101011100",
        2452 => "001101011010",
        2453 => "001101010111",
        2454 => "001101010101",
        2455 => "001101010010",
        2456 => "001101010000",
        2457 => "001101001101",
        2458 => "001101001010",
        2459 => "001101001000",
        2460 => "001101000101",
        2461 => "001101000011",
        2462 => "001101000000",
        2463 => "001100111110",
        2464 => "001100111011",
        2465 => "001100111001",
        2466 => "001100110110",
        2467 => "001100110100",
        2468 => "001100110001",
        2469 => "001100101111",
        2470 => "001100101100",
        2471 => "001100101010",
        2472 => "001100100111",
        2473 => "001100100101",
        2474 => "001100100010",
        2475 => "001100100000",
        2476 => "001100011101",
        2477 => "001100011011",
        2478 => "001100011000",
        2479 => "001100010110",
        2480 => "001100010011",
        2481 => "001100010001",
        2482 => "001100001110",
        2483 => "001100001100",
        2484 => "001100001001",
        2485 => "001100000111",
        2486 => "001100000101",
        2487 => "001100000010",
        2488 => "001100000000",
        2489 => "001011111101",
        2490 => "001011111011",
        2491 => "001011111000",
        2492 => "001011110110",
        2493 => "001011110011",
        2494 => "001011110001",
        2495 => "001011101111",
        2496 => "001011101100",
        2497 => "001011101010",
        2498 => "001011100111",
        2499 => "001011100101",
        2500 => "001011100010",
        2501 => "001011100000",
        2502 => "001011011110",
        2503 => "001011011011",
        2504 => "001011011001",
        2505 => "001011010110",
        2506 => "001011010100",
        2507 => "001011010010",
        2508 => "001011001111",
        2509 => "001011001101",
        2510 => "001011001010",
        2511 => "001011001000",
        2512 => "001011000110",
        2513 => "001011000011",
        2514 => "001011000001",
        2515 => "001010111111",
        2516 => "001010111100",
        2517 => "001010111010",
        2518 => "001010110111",
        2519 => "001010110101",
        2520 => "001010110011",
        2521 => "001010110000",
        2522 => "001010101110",
        2523 => "001010101100",
        2524 => "001010101001",
        2525 => "001010100111",
        2526 => "001010100101",
        2527 => "001010100010",
        2528 => "001010100000",
        2529 => "001010011110",
        2530 => "001010011011",
        2531 => "001010011001",
        2532 => "001010010111",
        2533 => "001010010100",
        2534 => "001010010010",
        2535 => "001010010000",
        2536 => "001010001101",
        2537 => "001010001011",
        2538 => "001010001001",
        2539 => "001010000111",
        2540 => "001010000100",
        2541 => "001010000010",
        2542 => "001010000000",
        2543 => "001001111101",
        2544 => "001001111011",
        2545 => "001001111001",
        2546 => "001001110111",
        2547 => "001001110100",
        2548 => "001001110010",
        2549 => "001001110000",
        2550 => "001001101110",
        2551 => "001001101011",
        2552 => "001001101001",
        2553 => "001001100111",
        2554 => "001001100101",
        2555 => "001001100010",
        2556 => "001001100000",
        2557 => "001001011110",
        2558 => "001001011100",
        2559 => "001001011001",
        2560 => "001001010111",
        2561 => "001001010101",
        2562 => "001001010011",
        2563 => "001001010001",
        2564 => "001001001110",
        2565 => "001001001100",
        2566 => "001001001010",
        2567 => "001001001000",
        2568 => "001001000110",
        2569 => "001001000011",
        2570 => "001001000001",
        2571 => "001000111111",
        2572 => "001000111101",
        2573 => "001000111011",
        2574 => "001000111000",
        2575 => "001000110110",
        2576 => "001000110100",
        2577 => "001000110010",
        2578 => "001000110000",
        2579 => "001000101110",
        2580 => "001000101011",
        2581 => "001000101001",
        2582 => "001000100111",
        2583 => "001000100101",
        2584 => "001000100011",
        2585 => "001000100001",
        2586 => "001000011111",
        2587 => "001000011100",
        2588 => "001000011010",
        2589 => "001000011000",
        2590 => "001000010110",
        2591 => "001000010100",
        2592 => "001000010010",
        2593 => "001000010000",
        2594 => "001000001110",
        2595 => "001000001100",
        2596 => "001000001001",
        2597 => "001000000111",
        2598 => "001000000101",
        2599 => "001000000011",
        2600 => "001000000001",
        2601 => "000111111111",
        2602 => "000111111101",
        2603 => "000111111011",
        2604 => "000111111001",
        2605 => "000111110111",
        2606 => "000111110101",
        2607 => "000111110011",
        2608 => "000111110001",
        2609 => "000111101111",
        2610 => "000111101101",
        2611 => "000111101010",
        2612 => "000111101000",
        2613 => "000111100110",
        2614 => "000111100100",
        2615 => "000111100010",
        2616 => "000111100000",
        2617 => "000111011110",
        2618 => "000111011100",
        2619 => "000111011010",
        2620 => "000111011000",
        2621 => "000111010110",
        2622 => "000111010100",
        2623 => "000111010010",
        2624 => "000111010000",
        2625 => "000111001110",
        2626 => "000111001100",
        2627 => "000111001010",
        2628 => "000111001000",
        2629 => "000111000110",
        2630 => "000111000100",
        2631 => "000111000010",
        2632 => "000111000000",
        2633 => "000110111110",
        2634 => "000110111101",
        2635 => "000110111011",
        2636 => "000110111001",
        2637 => "000110110111",
        2638 => "000110110101",
        2639 => "000110110011",
        2640 => "000110110001",
        2641 => "000110101111",
        2642 => "000110101101",
        2643 => "000110101011",
        2644 => "000110101001",
        2645 => "000110100111",
        2646 => "000110100101",
        2647 => "000110100011",
        2648 => "000110100010",
        2649 => "000110100000",
        2650 => "000110011110",
        2651 => "000110011100",
        2652 => "000110011010",
        2653 => "000110011000",
        2654 => "000110010110",
        2655 => "000110010100",
        2656 => "000110010010",
        2657 => "000110010001",
        2658 => "000110001111",
        2659 => "000110001101",
        2660 => "000110001011",
        2661 => "000110001001",
        2662 => "000110000111",
        2663 => "000110000101",
        2664 => "000110000100",
        2665 => "000110000010",
        2666 => "000110000000",
        2667 => "000101111110",
        2668 => "000101111100",
        2669 => "000101111010",
        2670 => "000101111001",
        2671 => "000101110111",
        2672 => "000101110101",
        2673 => "000101110011",
        2674 => "000101110001",
        2675 => "000101110000",
        2676 => "000101101110",
        2677 => "000101101100",
        2678 => "000101101010",
        2679 => "000101101000",
        2680 => "000101100111",
        2681 => "000101100101",
        2682 => "000101100011",
        2683 => "000101100001",
        2684 => "000101100000",
        2685 => "000101011110",
        2686 => "000101011100",
        2687 => "000101011010",
        2688 => "000101011001",
        2689 => "000101010111",
        2690 => "000101010101",
        2691 => "000101010011",
        2692 => "000101010010",
        2693 => "000101010000",
        2694 => "000101001110",
        2695 => "000101001100",
        2696 => "000101001011",
        2697 => "000101001001",
        2698 => "000101000111",
        2699 => "000101000110",
        2700 => "000101000100",
        2701 => "000101000010",
        2702 => "000101000001",
        2703 => "000100111111",
        2704 => "000100111101",
        2705 => "000100111011",
        2706 => "000100111010",
        2707 => "000100111000",
        2708 => "000100110110",
        2709 => "000100110101",
        2710 => "000100110011",
        2711 => "000100110001",
        2712 => "000100110000",
        2713 => "000100101110",
        2714 => "000100101101",
        2715 => "000100101011",
        2716 => "000100101001",
        2717 => "000100101000",
        2718 => "000100100110",
        2719 => "000100100100",
        2720 => "000100100011",
        2721 => "000100100001",
        2722 => "000100100000",
        2723 => "000100011110",
        2724 => "000100011100",
        2725 => "000100011011",
        2726 => "000100011001",
        2727 => "000100011000",
        2728 => "000100010110",
        2729 => "000100010100",
        2730 => "000100010011",
        2731 => "000100010001",
        2732 => "000100010000",
        2733 => "000100001110",
        2734 => "000100001101",
        2735 => "000100001011",
        2736 => "000100001001",
        2737 => "000100001000",
        2738 => "000100000110",
        2739 => "000100000101",
        2740 => "000100000011",
        2741 => "000100000010",
        2742 => "000100000000",
        2743 => "000011111111",
        2744 => "000011111101",
        2745 => "000011111100",
        2746 => "000011111010",
        2747 => "000011111001",
        2748 => "000011110111",
        2749 => "000011110110",
        2750 => "000011110100",
        2751 => "000011110011",
        2752 => "000011110001",
        2753 => "000011110000",
        2754 => "000011101110",
        2755 => "000011101101",
        2756 => "000011101011",
        2757 => "000011101010",
        2758 => "000011101000",
        2759 => "000011100111",
        2760 => "000011100110",
        2761 => "000011100100",
        2762 => "000011100011",
        2763 => "000011100001",
        2764 => "000011100000",
        2765 => "000011011110",
        2766 => "000011011101",
        2767 => "000011011100",
        2768 => "000011011010",
        2769 => "000011011001",
        2770 => "000011010111",
        2771 => "000011010110",
        2772 => "000011010101",
        2773 => "000011010011",
        2774 => "000011010010",
        2775 => "000011010000",
        2776 => "000011001111",
        2777 => "000011001110",
        2778 => "000011001100",
        2779 => "000011001011",
        2780 => "000011001001",
        2781 => "000011001000",
        2782 => "000011000111",
        2783 => "000011000101",
        2784 => "000011000100",
        2785 => "000011000011",
        2786 => "000011000001",
        2787 => "000011000000",
        2788 => "000010111111",
        2789 => "000010111101",
        2790 => "000010111100",
        2791 => "000010111011",
        2792 => "000010111001",
        2793 => "000010111000",
        2794 => "000010110111",
        2795 => "000010110110",
        2796 => "000010110100",
        2797 => "000010110011",
        2798 => "000010110010",
        2799 => "000010110000",
        2800 => "000010101111",
        2801 => "000010101110",
        2802 => "000010101101",
        2803 => "000010101011",
        2804 => "000010101010",
        2805 => "000010101001",
        2806 => "000010101000",
        2807 => "000010100110",
        2808 => "000010100101",
        2809 => "000010100100",
        2810 => "000010100011",
        2811 => "000010100001",
        2812 => "000010100000",
        2813 => "000010011111",
        2814 => "000010011110",
        2815 => "000010011101",
        2816 => "000010011011",
        2817 => "000010011010",
        2818 => "000010011001",
        2819 => "000010011000",
        2820 => "000010010111",
        2821 => "000010010101",
        2822 => "000010010100",
        2823 => "000010010011",
        2824 => "000010010010",
        2825 => "000010010001",
        2826 => "000010010000",
        2827 => "000010001110",
        2828 => "000010001101",
        2829 => "000010001100",
        2830 => "000010001011",
        2831 => "000010001010",
        2832 => "000010001001",
        2833 => "000010001000",
        2834 => "000010000110",
        2835 => "000010000101",
        2836 => "000010000100",
        2837 => "000010000011",
        2838 => "000010000010",
        2839 => "000010000001",
        2840 => "000010000000",
        2841 => "000001111111",
        2842 => "000001111110",
        2843 => "000001111101",
        2844 => "000001111011",
        2845 => "000001111010",
        2846 => "000001111001",
        2847 => "000001111000",
        2848 => "000001110111",
        2849 => "000001110110",
        2850 => "000001110101",
        2851 => "000001110100",
        2852 => "000001110011",
        2853 => "000001110010",
        2854 => "000001110001",
        2855 => "000001110000",
        2856 => "000001101111",
        2857 => "000001101110",
        2858 => "000001101101",
        2859 => "000001101100",
        2860 => "000001101011",
        2861 => "000001101010",
        2862 => "000001101001",
        2863 => "000001101000",
        2864 => "000001100111",
        2865 => "000001100110",
        2866 => "000001100101",
        2867 => "000001100100",
        2868 => "000001100011",
        2869 => "000001100010",
        2870 => "000001100001",
        2871 => "000001100000",
        2872 => "000001011111",
        2873 => "000001011110",
        2874 => "000001011101",
        2875 => "000001011100",
        2876 => "000001011011",
        2877 => "000001011010",
        2878 => "000001011001",
        2879 => "000001011001",
        2880 => "000001011000",
        2881 => "000001010111",
        2882 => "000001010110",
        2883 => "000001010101",
        2884 => "000001010100",
        2885 => "000001010011",
        2886 => "000001010010",
        2887 => "000001010001",
        2888 => "000001010001",
        2889 => "000001010000",
        2890 => "000001001111",
        2891 => "000001001110",
        2892 => "000001001101",
        2893 => "000001001100",
        2894 => "000001001011",
        2895 => "000001001011",
        2896 => "000001001010",
        2897 => "000001001001",
        2898 => "000001001000",
        2899 => "000001000111",
        2900 => "000001000110",
        2901 => "000001000110",
        2902 => "000001000101",
        2903 => "000001000100",
        2904 => "000001000011",
        2905 => "000001000010",
        2906 => "000001000010",
        2907 => "000001000001",
        2908 => "000001000000",
        2909 => "000000111111",
        2910 => "000000111110",
        2911 => "000000111110",
        2912 => "000000111101",
        2913 => "000000111100",
        2914 => "000000111011",
        2915 => "000000111011",
        2916 => "000000111010",
        2917 => "000000111001",
        2918 => "000000111000",
        2919 => "000000111000",
        2920 => "000000110111",
        2921 => "000000110110",
        2922 => "000000110101",
        2923 => "000000110101",
        2924 => "000000110100",
        2925 => "000000110011",
        2926 => "000000110011",
        2927 => "000000110010",
        2928 => "000000110001",
        2929 => "000000110001",
        2930 => "000000110000",
        2931 => "000000101111",
        2932 => "000000101111",
        2933 => "000000101110",
        2934 => "000000101101",
        2935 => "000000101101",
        2936 => "000000101100",
        2937 => "000000101011",
        2938 => "000000101011",
        2939 => "000000101010",
        2940 => "000000101001",
        2941 => "000000101001",
        2942 => "000000101000",
        2943 => "000000100111",
        2944 => "000000100111",
        2945 => "000000100110",
        2946 => "000000100110",
        2947 => "000000100101",
        2948 => "000000100100",
        2949 => "000000100100",
        2950 => "000000100011",
        2951 => "000000100011",
        2952 => "000000100010",
        2953 => "000000100010",
        2954 => "000000100001",
        2955 => "000000100000",
        2956 => "000000100000",
        2957 => "000000011111",
        2958 => "000000011111",
        2959 => "000000011110",
        2960 => "000000011110",
        2961 => "000000011101",
        2962 => "000000011101",
        2963 => "000000011100",
        2964 => "000000011100",
        2965 => "000000011011",
        2966 => "000000011011",
        2967 => "000000011010",
        2968 => "000000011010",
        2969 => "000000011001",
        2970 => "000000011001",
        2971 => "000000011000",
        2972 => "000000011000",
        2973 => "000000010111",
        2974 => "000000010111",
        2975 => "000000010110",
        2976 => "000000010110",
        2977 => "000000010101",
        2978 => "000000010101",
        2979 => "000000010100",
        2980 => "000000010100",
        2981 => "000000010011",
        2982 => "000000010011",
        2983 => "000000010011",
        2984 => "000000010010",
        2985 => "000000010010",
        2986 => "000000010001",
        2987 => "000000010001",
        2988 => "000000010000",
        2989 => "000000010000",
        2990 => "000000010000",
        2991 => "000000001111",
        2992 => "000000001111",
        2993 => "000000001111",
        2994 => "000000001110",
        2995 => "000000001110",
        2996 => "000000001101",
        2997 => "000000001101",
        2998 => "000000001101",
        2999 => "000000001100",
        3000 => "000000001100",
        3001 => "000000001100",
        3002 => "000000001011",
        3003 => "000000001011",
        3004 => "000000001011",
        3005 => "000000001010",
        3006 => "000000001010",
        3007 => "000000001010",
        3008 => "000000001001",
        3009 => "000000001001",
        3010 => "000000001001",
        3011 => "000000001000",
        3012 => "000000001000",
        3013 => "000000001000",
        3014 => "000000001000",
        3015 => "000000000111",
        3016 => "000000000111",
        3017 => "000000000111",
        3018 => "000000000111",
        3019 => "000000000110",
        3020 => "000000000110",
        3021 => "000000000110",
        3022 => "000000000110",
        3023 => "000000000101",
        3024 => "000000000101",
        3025 => "000000000101",
        3026 => "000000000101",
        3027 => "000000000100",
        3028 => "000000000100",
        3029 => "000000000100",
        3030 => "000000000100",
        3031 => "000000000100",
        3032 => "000000000011",
        3033 => "000000000011",
        3034 => "000000000011",
        3035 => "000000000011",
        3036 => "000000000011",
        3037 => "000000000010",
        3038 => "000000000010",
        3039 => "000000000010",
        3040 => "000000000010",
        3041 => "000000000010",
        3042 => "000000000010",
        3043 => "000000000010",
        3044 => "000000000001",
        3045 => "000000000001",
        3046 => "000000000001",
        3047 => "000000000001",
        3048 => "000000000001",
        3049 => "000000000001",
        3050 => "000000000001",
        3051 => "000000000001",
        3052 => "000000000000",
        3053 => "000000000000",
        3054 => "000000000000",
        3055 => "000000000000",
        3056 => "000000000000",
        3057 => "000000000000",
        3058 => "000000000000",
        3059 => "000000000000",
        3060 => "000000000000",
        3061 => "000000000000",
        3062 => "000000000000",
        3063 => "000000000000",
        3064 => "000000000000",
        3065 => "000000000000",
        3066 => "000000000000",
        3067 => "000000000000",
        3068 => "000000000000",
        3069 => "000000000000",
        3070 => "000000000000",
        3071 => "000000000000",
        3072 => "000000000000",
        3073 => "000000000000",
        3074 => "000000000000",
        3075 => "000000000000",
        3076 => "000000000000",
        3077 => "000000000000",
        3078 => "000000000000",
        3079 => "000000000000",
        3080 => "000000000000",
        3081 => "000000000000",
        3082 => "000000000000",
        3083 => "000000000000",
        3084 => "000000000000",
        3085 => "000000000000",
        3086 => "000000000000",
        3087 => "000000000000",
        3088 => "000000000000",
        3089 => "000000000000",
        3090 => "000000000000",
        3091 => "000000000000",
        3092 => "000000000000",
        3093 => "000000000001",
        3094 => "000000000001",
        3095 => "000000000001",
        3096 => "000000000001",
        3097 => "000000000001",
        3098 => "000000000001",
        3099 => "000000000001",
        3100 => "000000000001",
        3101 => "000000000010",
        3102 => "000000000010",
        3103 => "000000000010",
        3104 => "000000000010",
        3105 => "000000000010",
        3106 => "000000000010",
        3107 => "000000000010",
        3108 => "000000000011",
        3109 => "000000000011",
        3110 => "000000000011",
        3111 => "000000000011",
        3112 => "000000000011",
        3113 => "000000000100",
        3114 => "000000000100",
        3115 => "000000000100",
        3116 => "000000000100",
        3117 => "000000000100",
        3118 => "000000000101",
        3119 => "000000000101",
        3120 => "000000000101",
        3121 => "000000000101",
        3122 => "000000000110",
        3123 => "000000000110",
        3124 => "000000000110",
        3125 => "000000000110",
        3126 => "000000000111",
        3127 => "000000000111",
        3128 => "000000000111",
        3129 => "000000000111",
        3130 => "000000001000",
        3131 => "000000001000",
        3132 => "000000001000",
        3133 => "000000001000",
        3134 => "000000001001",
        3135 => "000000001001",
        3136 => "000000001001",
        3137 => "000000001010",
        3138 => "000000001010",
        3139 => "000000001010",
        3140 => "000000001011",
        3141 => "000000001011",
        3142 => "000000001011",
        3143 => "000000001100",
        3144 => "000000001100",
        3145 => "000000001100",
        3146 => "000000001101",
        3147 => "000000001101",
        3148 => "000000001101",
        3149 => "000000001110",
        3150 => "000000001110",
        3151 => "000000001111",
        3152 => "000000001111",
        3153 => "000000001111",
        3154 => "000000010000",
        3155 => "000000010000",
        3156 => "000000010000",
        3157 => "000000010001",
        3158 => "000000010001",
        3159 => "000000010010",
        3160 => "000000010010",
        3161 => "000000010011",
        3162 => "000000010011",
        3163 => "000000010011",
        3164 => "000000010100",
        3165 => "000000010100",
        3166 => "000000010101",
        3167 => "000000010101",
        3168 => "000000010110",
        3169 => "000000010110",
        3170 => "000000010111",
        3171 => "000000010111",
        3172 => "000000011000",
        3173 => "000000011000",
        3174 => "000000011001",
        3175 => "000000011001",
        3176 => "000000011010",
        3177 => "000000011010",
        3178 => "000000011011",
        3179 => "000000011011",
        3180 => "000000011100",
        3181 => "000000011100",
        3182 => "000000011101",
        3183 => "000000011101",
        3184 => "000000011110",
        3185 => "000000011110",
        3186 => "000000011111",
        3187 => "000000011111",
        3188 => "000000100000",
        3189 => "000000100000",
        3190 => "000000100001",
        3191 => "000000100010",
        3192 => "000000100010",
        3193 => "000000100011",
        3194 => "000000100011",
        3195 => "000000100100",
        3196 => "000000100100",
        3197 => "000000100101",
        3198 => "000000100110",
        3199 => "000000100110",
        3200 => "000000100111",
        3201 => "000000100111",
        3202 => "000000101000",
        3203 => "000000101001",
        3204 => "000000101001",
        3205 => "000000101010",
        3206 => "000000101011",
        3207 => "000000101011",
        3208 => "000000101100",
        3209 => "000000101101",
        3210 => "000000101101",
        3211 => "000000101110",
        3212 => "000000101111",
        3213 => "000000101111",
        3214 => "000000110000",
        3215 => "000000110001",
        3216 => "000000110001",
        3217 => "000000110010",
        3218 => "000000110011",
        3219 => "000000110011",
        3220 => "000000110100",
        3221 => "000000110101",
        3222 => "000000110101",
        3223 => "000000110110",
        3224 => "000000110111",
        3225 => "000000111000",
        3226 => "000000111000",
        3227 => "000000111001",
        3228 => "000000111010",
        3229 => "000000111011",
        3230 => "000000111011",
        3231 => "000000111100",
        3232 => "000000111101",
        3233 => "000000111110",
        3234 => "000000111110",
        3235 => "000000111111",
        3236 => "000001000000",
        3237 => "000001000001",
        3238 => "000001000010",
        3239 => "000001000010",
        3240 => "000001000011",
        3241 => "000001000100",
        3242 => "000001000101",
        3243 => "000001000110",
        3244 => "000001000110",
        3245 => "000001000111",
        3246 => "000001001000",
        3247 => "000001001001",
        3248 => "000001001010",
        3249 => "000001001011",
        3250 => "000001001011",
        3251 => "000001001100",
        3252 => "000001001101",
        3253 => "000001001110",
        3254 => "000001001111",
        3255 => "000001010000",
        3256 => "000001010001",
        3257 => "000001010001",
        3258 => "000001010010",
        3259 => "000001010011",
        3260 => "000001010100",
        3261 => "000001010101",
        3262 => "000001010110",
        3263 => "000001010111",
        3264 => "000001011000",
        3265 => "000001011001",
        3266 => "000001011001",
        3267 => "000001011010",
        3268 => "000001011011",
        3269 => "000001011100",
        3270 => "000001011101",
        3271 => "000001011110",
        3272 => "000001011111",
        3273 => "000001100000",
        3274 => "000001100001",
        3275 => "000001100010",
        3276 => "000001100011",
        3277 => "000001100100",
        3278 => "000001100101",
        3279 => "000001100110",
        3280 => "000001100111",
        3281 => "000001101000",
        3282 => "000001101001",
        3283 => "000001101010",
        3284 => "000001101011",
        3285 => "000001101100",
        3286 => "000001101101",
        3287 => "000001101110",
        3288 => "000001101111",
        3289 => "000001110000",
        3290 => "000001110001",
        3291 => "000001110010",
        3292 => "000001110011",
        3293 => "000001110100",
        3294 => "000001110101",
        3295 => "000001110110",
        3296 => "000001110111",
        3297 => "000001111000",
        3298 => "000001111001",
        3299 => "000001111010",
        3300 => "000001111011",
        3301 => "000001111101",
        3302 => "000001111110",
        3303 => "000001111111",
        3304 => "000010000000",
        3305 => "000010000001",
        3306 => "000010000010",
        3307 => "000010000011",
        3308 => "000010000100",
        3309 => "000010000101",
        3310 => "000010000110",
        3311 => "000010001000",
        3312 => "000010001001",
        3313 => "000010001010",
        3314 => "000010001011",
        3315 => "000010001100",
        3316 => "000010001101",
        3317 => "000010001110",
        3318 => "000010010000",
        3319 => "000010010001",
        3320 => "000010010010",
        3321 => "000010010011",
        3322 => "000010010100",
        3323 => "000010010101",
        3324 => "000010010111",
        3325 => "000010011000",
        3326 => "000010011001",
        3327 => "000010011010",
        3328 => "000010011011",
        3329 => "000010011101",
        3330 => "000010011110",
        3331 => "000010011111",
        3332 => "000010100000",
        3333 => "000010100001",
        3334 => "000010100011",
        3335 => "000010100100",
        3336 => "000010100101",
        3337 => "000010100110",
        3338 => "000010101000",
        3339 => "000010101001",
        3340 => "000010101010",
        3341 => "000010101011",
        3342 => "000010101101",
        3343 => "000010101110",
        3344 => "000010101111",
        3345 => "000010110000",
        3346 => "000010110010",
        3347 => "000010110011",
        3348 => "000010110100",
        3349 => "000010110110",
        3350 => "000010110111",
        3351 => "000010111000",
        3352 => "000010111001",
        3353 => "000010111011",
        3354 => "000010111100",
        3355 => "000010111101",
        3356 => "000010111111",
        3357 => "000011000000",
        3358 => "000011000001",
        3359 => "000011000011",
        3360 => "000011000100",
        3361 => "000011000101",
        3362 => "000011000111",
        3363 => "000011001000",
        3364 => "000011001001",
        3365 => "000011001011",
        3366 => "000011001100",
        3367 => "000011001110",
        3368 => "000011001111",
        3369 => "000011010000",
        3370 => "000011010010",
        3371 => "000011010011",
        3372 => "000011010101",
        3373 => "000011010110",
        3374 => "000011010111",
        3375 => "000011011001",
        3376 => "000011011010",
        3377 => "000011011100",
        3378 => "000011011101",
        3379 => "000011011110",
        3380 => "000011100000",
        3381 => "000011100001",
        3382 => "000011100011",
        3383 => "000011100100",
        3384 => "000011100110",
        3385 => "000011100111",
        3386 => "000011101000",
        3387 => "000011101010",
        3388 => "000011101011",
        3389 => "000011101101",
        3390 => "000011101110",
        3391 => "000011110000",
        3392 => "000011110001",
        3393 => "000011110011",
        3394 => "000011110100",
        3395 => "000011110110",
        3396 => "000011110111",
        3397 => "000011111001",
        3398 => "000011111010",
        3399 => "000011111100",
        3400 => "000011111101",
        3401 => "000011111111",
        3402 => "000100000000",
        3403 => "000100000010",
        3404 => "000100000011",
        3405 => "000100000101",
        3406 => "000100000110",
        3407 => "000100001000",
        3408 => "000100001001",
        3409 => "000100001011",
        3410 => "000100001101",
        3411 => "000100001110",
        3412 => "000100010000",
        3413 => "000100010001",
        3414 => "000100010011",
        3415 => "000100010100",
        3416 => "000100010110",
        3417 => "000100011000",
        3418 => "000100011001",
        3419 => "000100011011",
        3420 => "000100011100",
        3421 => "000100011110",
        3422 => "000100100000",
        3423 => "000100100001",
        3424 => "000100100011",
        3425 => "000100100100",
        3426 => "000100100110",
        3427 => "000100101000",
        3428 => "000100101001",
        3429 => "000100101011",
        3430 => "000100101101",
        3431 => "000100101110",
        3432 => "000100110000",
        3433 => "000100110001",
        3434 => "000100110011",
        3435 => "000100110101",
        3436 => "000100110110",
        3437 => "000100111000",
        3438 => "000100111010",
        3439 => "000100111011",
        3440 => "000100111101",
        3441 => "000100111111",
        3442 => "000101000001",
        3443 => "000101000010",
        3444 => "000101000100",
        3445 => "000101000110",
        3446 => "000101000111",
        3447 => "000101001001",
        3448 => "000101001011",
        3449 => "000101001100",
        3450 => "000101001110",
        3451 => "000101010000",
        3452 => "000101010010",
        3453 => "000101010011",
        3454 => "000101010101",
        3455 => "000101010111",
        3456 => "000101011001",
        3457 => "000101011010",
        3458 => "000101011100",
        3459 => "000101011110",
        3460 => "000101100000",
        3461 => "000101100001",
        3462 => "000101100011",
        3463 => "000101100101",
        3464 => "000101100111",
        3465 => "000101101000",
        3466 => "000101101010",
        3467 => "000101101100",
        3468 => "000101101110",
        3469 => "000101110000",
        3470 => "000101110001",
        3471 => "000101110011",
        3472 => "000101110101",
        3473 => "000101110111",
        3474 => "000101111001",
        3475 => "000101111010",
        3476 => "000101111100",
        3477 => "000101111110",
        3478 => "000110000000",
        3479 => "000110000010",
        3480 => "000110000100",
        3481 => "000110000101",
        3482 => "000110000111",
        3483 => "000110001001",
        3484 => "000110001011",
        3485 => "000110001101",
        3486 => "000110001111",
        3487 => "000110010001",
        3488 => "000110010010",
        3489 => "000110010100",
        3490 => "000110010110",
        3491 => "000110011000",
        3492 => "000110011010",
        3493 => "000110011100",
        3494 => "000110011110",
        3495 => "000110100000",
        3496 => "000110100010",
        3497 => "000110100011",
        3498 => "000110100101",
        3499 => "000110100111",
        3500 => "000110101001",
        3501 => "000110101011",
        3502 => "000110101101",
        3503 => "000110101111",
        3504 => "000110110001",
        3505 => "000110110011",
        3506 => "000110110101",
        3507 => "000110110111",
        3508 => "000110111001",
        3509 => "000110111011",
        3510 => "000110111101",
        3511 => "000110111110",
        3512 => "000111000000",
        3513 => "000111000010",
        3514 => "000111000100",
        3515 => "000111000110",
        3516 => "000111001000",
        3517 => "000111001010",
        3518 => "000111001100",
        3519 => "000111001110",
        3520 => "000111010000",
        3521 => "000111010010",
        3522 => "000111010100",
        3523 => "000111010110",
        3524 => "000111011000",
        3525 => "000111011010",
        3526 => "000111011100",
        3527 => "000111011110",
        3528 => "000111100000",
        3529 => "000111100010",
        3530 => "000111100100",
        3531 => "000111100110",
        3532 => "000111101000",
        3533 => "000111101010",
        3534 => "000111101101",
        3535 => "000111101111",
        3536 => "000111110001",
        3537 => "000111110011",
        3538 => "000111110101",
        3539 => "000111110111",
        3540 => "000111111001",
        3541 => "000111111011",
        3542 => "000111111101",
        3543 => "000111111111",
        3544 => "001000000001",
        3545 => "001000000011",
        3546 => "001000000101",
        3547 => "001000000111",
        3548 => "001000001001",
        3549 => "001000001100",
        3550 => "001000001110",
        3551 => "001000010000",
        3552 => "001000010010",
        3553 => "001000010100",
        3554 => "001000010110",
        3555 => "001000011000",
        3556 => "001000011010",
        3557 => "001000011100",
        3558 => "001000011111",
        3559 => "001000100001",
        3560 => "001000100011",
        3561 => "001000100101",
        3562 => "001000100111",
        3563 => "001000101001",
        3564 => "001000101011",
        3565 => "001000101110",
        3566 => "001000110000",
        3567 => "001000110010",
        3568 => "001000110100",
        3569 => "001000110110",
        3570 => "001000111000",
        3571 => "001000111011",
        3572 => "001000111101",
        3573 => "001000111111",
        3574 => "001001000001",
        3575 => "001001000011",
        3576 => "001001000110",
        3577 => "001001001000",
        3578 => "001001001010",
        3579 => "001001001100",
        3580 => "001001001110",
        3581 => "001001010001",
        3582 => "001001010011",
        3583 => "001001010101",
        3584 => "001001010111",
        3585 => "001001011001",
        3586 => "001001011100",
        3587 => "001001011110",
        3588 => "001001100000",
        3589 => "001001100010",
        3590 => "001001100101",
        3591 => "001001100111",
        3592 => "001001101001",
        3593 => "001001101011",
        3594 => "001001101110",
        3595 => "001001110000",
        3596 => "001001110010",
        3597 => "001001110100",
        3598 => "001001110111",
        3599 => "001001111001",
        3600 => "001001111011",
        3601 => "001001111101",
        3602 => "001010000000",
        3603 => "001010000010",
        3604 => "001010000100",
        3605 => "001010000111",
        3606 => "001010001001",
        3607 => "001010001011",
        3608 => "001010001101",
        3609 => "001010010000",
        3610 => "001010010010",
        3611 => "001010010100",
        3612 => "001010010111",
        3613 => "001010011001",
        3614 => "001010011011",
        3615 => "001010011110",
        3616 => "001010100000",
        3617 => "001010100010",
        3618 => "001010100101",
        3619 => "001010100111",
        3620 => "001010101001",
        3621 => "001010101100",
        3622 => "001010101110",
        3623 => "001010110000",
        3624 => "001010110011",
        3625 => "001010110101",
        3626 => "001010110111",
        3627 => "001010111010",
        3628 => "001010111100",
        3629 => "001010111111",
        3630 => "001011000001",
        3631 => "001011000011",
        3632 => "001011000110",
        3633 => "001011001000",
        3634 => "001011001010",
        3635 => "001011001101",
        3636 => "001011001111",
        3637 => "001011010010",
        3638 => "001011010100",
        3639 => "001011010110",
        3640 => "001011011001",
        3641 => "001011011011",
        3642 => "001011011110",
        3643 => "001011100000",
        3644 => "001011100010",
        3645 => "001011100101",
        3646 => "001011100111",
        3647 => "001011101010",
        3648 => "001011101100",
        3649 => "001011101111",
        3650 => "001011110001",
        3651 => "001011110011",
        3652 => "001011110110",
        3653 => "001011111000",
        3654 => "001011111011",
        3655 => "001011111101",
        3656 => "001100000000",
        3657 => "001100000010",
        3658 => "001100000101",
        3659 => "001100000111",
        3660 => "001100001001",
        3661 => "001100001100",
        3662 => "001100001110",
        3663 => "001100010001",
        3664 => "001100010011",
        3665 => "001100010110",
        3666 => "001100011000",
        3667 => "001100011011",
        3668 => "001100011101",
        3669 => "001100100000",
        3670 => "001100100010",
        3671 => "001100100101",
        3672 => "001100100111",
        3673 => "001100101010",
        3674 => "001100101100",
        3675 => "001100101111",
        3676 => "001100110001",
        3677 => "001100110100",
        3678 => "001100110110",
        3679 => "001100111001",
        3680 => "001100111011",
        3681 => "001100111110",
        3682 => "001101000000",
        3683 => "001101000011",
        3684 => "001101000101",
        3685 => "001101001000",
        3686 => "001101001010",
        3687 => "001101001101",
        3688 => "001101010000",
        3689 => "001101010010",
        3690 => "001101010101",
        3691 => "001101010111",
        3692 => "001101011010",
        3693 => "001101011100",
        3694 => "001101011111",
        3695 => "001101100001",
        3696 => "001101100100",
        3697 => "001101100111",
        3698 => "001101101001",
        3699 => "001101101100",
        3700 => "001101101110",
        3701 => "001101110001",
        3702 => "001101110011",
        3703 => "001101110110",
        3704 => "001101111001",
        3705 => "001101111011",
        3706 => "001101111110",
        3707 => "001110000000",
        3708 => "001110000011",
        3709 => "001110000110",
        3710 => "001110001000",
        3711 => "001110001011",
        3712 => "001110001101",
        3713 => "001110010000",
        3714 => "001110010011",
        3715 => "001110010101",
        3716 => "001110011000",
        3717 => "001110011011",
        3718 => "001110011101",
        3719 => "001110100000",
        3720 => "001110100010",
        3721 => "001110100101",
        3722 => "001110101000",
        3723 => "001110101010",
        3724 => "001110101101",
        3725 => "001110110000",
        3726 => "001110110010",
        3727 => "001110110101",
        3728 => "001110111000",
        3729 => "001110111010",
        3730 => "001110111101",
        3731 => "001111000000",
        3732 => "001111000010",
        3733 => "001111000101",
        3734 => "001111001000",
        3735 => "001111001010",
        3736 => "001111001101",
        3737 => "001111010000",
        3738 => "001111010010",
        3739 => "001111010101",
        3740 => "001111011000",
        3741 => "001111011010",
        3742 => "001111011101",
        3743 => "001111100000",
        3744 => "001111100010",
        3745 => "001111100101",
        3746 => "001111101000",
        3747 => "001111101010",
        3748 => "001111101101",
        3749 => "001111110000",
        3750 => "001111110011",
        3751 => "001111110101",
        3752 => "001111111000",
        3753 => "001111111011",
        3754 => "001111111101",
        3755 => "010000000000",
        3756 => "010000000011",
        3757 => "010000000110",
        3758 => "010000001000",
        3759 => "010000001011",
        3760 => "010000001110",
        3761 => "010000010001",
        3762 => "010000010011",
        3763 => "010000010110",
        3764 => "010000011001",
        3765 => "010000011011",
        3766 => "010000011110",
        3767 => "010000100001",
        3768 => "010000100100",
        3769 => "010000100110",
        3770 => "010000101001",
        3771 => "010000101100",
        3772 => "010000101111",
        3773 => "010000110010",
        3774 => "010000110100",
        3775 => "010000110111",
        3776 => "010000111010",
        3777 => "010000111101",
        3778 => "010000111111",
        3779 => "010001000010",
        3780 => "010001000101",
        3781 => "010001001000",
        3782 => "010001001010",
        3783 => "010001001101",
        3784 => "010001010000",
        3785 => "010001010011",
        3786 => "010001010110",
        3787 => "010001011000",
        3788 => "010001011011",
        3789 => "010001011110",
        3790 => "010001100001",
        3791 => "010001100100",
        3792 => "010001100110",
        3793 => "010001101001",
        3794 => "010001101100",
        3795 => "010001101111",
        3796 => "010001110010",
        3797 => "010001110100",
        3798 => "010001110111",
        3799 => "010001111010",
        3800 => "010001111101",
        3801 => "010010000000",
        3802 => "010010000011",
        3803 => "010010000101",
        3804 => "010010001000",
        3805 => "010010001011",
        3806 => "010010001110",
        3807 => "010010010001",
        3808 => "010010010100",
        3809 => "010010010110",
        3810 => "010010011001",
        3811 => "010010011100",
        3812 => "010010011111",
        3813 => "010010100010",
        3814 => "010010100101",
        3815 => "010010101000",
        3816 => "010010101010",
        3817 => "010010101101",
        3818 => "010010110000",
        3819 => "010010110011",
        3820 => "010010110110",
        3821 => "010010111001",
        3822 => "010010111100",
        3823 => "010010111110",
        3824 => "010011000001",
        3825 => "010011000100",
        3826 => "010011000111",
        3827 => "010011001010",
        3828 => "010011001101",
        3829 => "010011010000",
        3830 => "010011010011",
        3831 => "010011010101",
        3832 => "010011011000",
        3833 => "010011011011",
        3834 => "010011011110",
        3835 => "010011100001",
        3836 => "010011100100",
        3837 => "010011100111",
        3838 => "010011101010",
        3839 => "010011101101",
        3840 => "010011101111",
        3841 => "010011110010",
        3842 => "010011110101",
        3843 => "010011111000",
        3844 => "010011111011",
        3845 => "010011111110",
        3846 => "010100000001",
        3847 => "010100000100",
        3848 => "010100000111",
        3849 => "010100001010",
        3850 => "010100001101",
        3851 => "010100001111",
        3852 => "010100010010",
        3853 => "010100010101",
        3854 => "010100011000",
        3855 => "010100011011",
        3856 => "010100011110",
        3857 => "010100100001",
        3858 => "010100100100",
        3859 => "010100100111",
        3860 => "010100101010",
        3861 => "010100101101",
        3862 => "010100110000",
        3863 => "010100110011",
        3864 => "010100110110",
        3865 => "010100111001",
        3866 => "010100111100",
        3867 => "010100111110",
        3868 => "010101000001",
        3869 => "010101000100",
        3870 => "010101000111",
        3871 => "010101001010",
        3872 => "010101001101",
        3873 => "010101010000",
        3874 => "010101010011",
        3875 => "010101010110",
        3876 => "010101011001",
        3877 => "010101011100",
        3878 => "010101011111",
        3879 => "010101100010",
        3880 => "010101100101",
        3881 => "010101101000",
        3882 => "010101101011",
        3883 => "010101101110",
        3884 => "010101110001",
        3885 => "010101110100",
        3886 => "010101110111",
        3887 => "010101111010",
        3888 => "010101111101",
        3889 => "010110000000",
        3890 => "010110000011",
        3891 => "010110000110",
        3892 => "010110001001",
        3893 => "010110001100",
        3894 => "010110001111",
        3895 => "010110010010",
        3896 => "010110010101",
        3897 => "010110011000",
        3898 => "010110011011",
        3899 => "010110011110",
        3900 => "010110100001",
        3901 => "010110100100",
        3902 => "010110100111",
        3903 => "010110101010",
        3904 => "010110101101",
        3905 => "010110110000",
        3906 => "010110110011",
        3907 => "010110110110",
        3908 => "010110111001",
        3909 => "010110111100",
        3910 => "010110111111",
        3911 => "010111000010",
        3912 => "010111000101",
        3913 => "010111001000",
        3914 => "010111001011",
        3915 => "010111001110",
        3916 => "010111010001",
        3917 => "010111010100",
        3918 => "010111010111",
        3919 => "010111011010",
        3920 => "010111011101",
        3921 => "010111100000",
        3922 => "010111100011",
        3923 => "010111100110",
        3924 => "010111101001",
        3925 => "010111101100",
        3926 => "010111101111",
        3927 => "010111110010",
        3928 => "010111110101",
        3929 => "010111111000",
        3930 => "010111111011",
        3931 => "010111111110",
        3932 => "011000000001",
        3933 => "011000000100",
        3934 => "011000000111",
        3935 => "011000001010",
        3936 => "011000001101",
        3937 => "011000010001",
        3938 => "011000010100",
        3939 => "011000010111",
        3940 => "011000011010",
        3941 => "011000011101",
        3942 => "011000100000",
        3943 => "011000100011",
        3944 => "011000100110",
        3945 => "011000101001",
        3946 => "011000101100",
        3947 => "011000101111",
        3948 => "011000110010",
        3949 => "011000110101",
        3950 => "011000111000",
        3951 => "011000111011",
        3952 => "011000111110",
        3953 => "011001000001",
        3954 => "011001000101",
        3955 => "011001001000",
        3956 => "011001001011",
        3957 => "011001001110",
        3958 => "011001010001",
        3959 => "011001010100",
        3960 => "011001010111",
        3961 => "011001011010",
        3962 => "011001011101",
        3963 => "011001100000",
        3964 => "011001100011",
        3965 => "011001100110",
        3966 => "011001101001",
        3967 => "011001101100",
        3968 => "011001110000",
        3969 => "011001110011",
        3970 => "011001110110",
        3971 => "011001111001",
        3972 => "011001111100",
        3973 => "011001111111",
        3974 => "011010000010",
        3975 => "011010000101",
        3976 => "011010001000",
        3977 => "011010001011",
        3978 => "011010001110",
        3979 => "011010010001",
        3980 => "011010010101",
        3981 => "011010011000",
        3982 => "011010011011",
        3983 => "011010011110",
        3984 => "011010100001",
        3985 => "011010100100",
        3986 => "011010100111",
        3987 => "011010101010",
        3988 => "011010101101",
        3989 => "011010110000",
        3990 => "011010110100",
        3991 => "011010110111",
        3992 => "011010111010",
        3993 => "011010111101",
        3994 => "011011000000",
        3995 => "011011000011",
        3996 => "011011000110",
        3997 => "011011001001",
        3998 => "011011001100",
        3999 => "011011001111",
        4000 => "011011010011",
        4001 => "011011010110",
        4002 => "011011011001",
        4003 => "011011011100",
        4004 => "011011011111",
        4005 => "011011100010",
        4006 => "011011100101",
        4007 => "011011101000",
        4008 => "011011101011",
        4009 => "011011101111",
        4010 => "011011110010",
        4011 => "011011110101",
        4012 => "011011111000",
        4013 => "011011111011",
        4014 => "011011111110",
        4015 => "011100000001",
        4016 => "011100000100",
        4017 => "011100000111",
        4018 => "011100001011",
        4019 => "011100001110",
        4020 => "011100010001",
        4021 => "011100010100",
        4022 => "011100010111",
        4023 => "011100011010",
        4024 => "011100011101",
        4025 => "011100100000",
        4026 => "011100100100",
        4027 => "011100100111",
        4028 => "011100101010",
        4029 => "011100101101",
        4030 => "011100110000",
        4031 => "011100110011",
        4032 => "011100110110",
        4033 => "011100111001",
        4034 => "011100111101",
        4035 => "011101000000",
        4036 => "011101000011",
        4037 => "011101000110",
        4038 => "011101001001",
        4039 => "011101001100",
        4040 => "011101001111",
        4041 => "011101010010",
        4042 => "011101010110",
        4043 => "011101011001",
        4044 => "011101011100",
        4045 => "011101011111",
        4046 => "011101100010",
        4047 => "011101100101",
        4048 => "011101101000",
        4049 => "011101101100",
        4050 => "011101101111",
        4051 => "011101110010",
        4052 => "011101110101",
        4053 => "011101111000",
        4054 => "011101111011",
        4055 => "011101111110",
        4056 => "011110000001",
        4057 => "011110000101",
        4058 => "011110001000",
        4059 => "011110001011",
        4060 => "011110001110",
        4061 => "011110010001",
        4062 => "011110010100",
        4063 => "011110010111",
        4064 => "011110011011",
        4065 => "011110011110",
        4066 => "011110100001",
        4067 => "011110100100",
        4068 => "011110100111",
        4069 => "011110101010",
        4070 => "011110101101",
        4071 => "011110110000",
        4072 => "011110110100",
        4073 => "011110110111",
        4074 => "011110111010",
        4075 => "011110111101",
        4076 => "011111000000",
        4077 => "011111000011",
        4078 => "011111000110",
        4079 => "011111001010",
        4080 => "011111001101",
        4081 => "011111010000",
        4082 => "011111010011",
        4083 => "011111010110",
        4084 => "011111011001",
        4085 => "011111011100",
        4086 => "011111100000",
        4087 => "011111100011",
        4088 => "011111100110",
        4089 => "011111101001",
        4090 => "011111101100",
        4091 => "011111101111",
        4092 => "011111110010",
        4093 => "011111110110",
        4094 => "011111111001",
        4095 => "011111111100");

    signal phase_accum: std_logic_vector(15 downto 0);
    signal lut_value: std_logic_vector(11 downto 0);
    signal probe_out: std_logic_vector(11 downto 0);
    signal probe_pha: std_logic_vector(15 downto 0);

begin
        -- behavior
    process(clk_i)
        begin 
            if rising_edge(clk_i) then
                if rst_i = '1' then
                    phase_accum <= (others => '0');
                else 
                    phase_accum <= std_logic_vector(unsigned(phase_accum) + unsigned(probe_pha));
            end if;
        end if; 
        end process;

        lut_value <= std_logic_vector(unsigned(phase_accum(15 downto 4)));

    probe_out <= sin_lut(to_integer(unsigned(lut_value)));
    
    ila_inst : ila_0
    PORT MAP (
        clk => clk_i,
        probe0 => probe_out
    );
    
    vio_inst : vio_0
      PORT MAP (
        clk => clk_i,
        probe_out0 => probe_pha
      );

end architecture;